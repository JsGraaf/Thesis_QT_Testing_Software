

module lut_2_ro(
   input en,
   output out,
);

(*keep*)wire connect;

assign connect = en ? connect : 0;
assign out = en ? connect : 0;

LUT2 #(
   .INIT(4'b0001)
) ro (
   .I0(connect),
   .I1(1'b0),
   .O(out)
);
endmodule

 
module eightbitadd ( 
      input wire [31:0] a,
      input wire [31:0] b,
      input c_in,
      output reg c_out,
      output reg[31:0] sum,
      input clk,);

   always @ (posedge clk) begin
      {c_out, sum} = a + b + c_in;
   end
endmodule

module doubleeightbitadd (
   input wire [31:0] a1,
   input wire [31:0] a2,
   input wire [31:0] b1,
   input wire [31:0] b2,
   output wire [31:0] sum,
   input clk,);

wire [31:0] sum1;
wire [31:0] sum2;

 eightbitadd add1(
   .a(a1),
   .b(a2),
   .c_in(1'b0),
   .sum(sum1),
   .clk(clk),
);

 eightbitadd add2(
   .a(b1),
   .b(b2),
   .c_in(1'b0),
   .sum(sum2),
   .clk(clk),
);

 eightbitadd addTot(
   .a(sum1),
   .b(sum2),
   .c_in(1'b0),
   .sum(sum),
   .clk(clk),
);
endmodule

module quadeightbitadd (
   input wire [31:0] a1,
   input wire [31:0] a2,
   input wire [31:0] a3,
   input wire [31:0] a4,
   input wire [31:0] b1,
   input wire [31:0] b2,
   input wire [31:0] b3,
   input wire [31:0] b4,
   output wire[31:0] sum,
   input clk,
);

reg [31:0] sum1;
reg [31:0] sum2;

doubleeightbitadd add1(
   .a1(a1),
   .a2(a2),
   .b1(a3),
   .b2(a4),
   .clk(clk),
   .sum(sum1),
);

doubleeightbitadd add2(
   .a1(b1),
   .a2(b2),
   .b1(b3),
   .b2(b4),
   .clk(clk),
   .sum(sum2),
);

eightbitadd addTot(
   .a(sum1),
   .b(sum2),
   .c_in(1'b0),
   .clk(clk),
   .sum(sum),
);
endmodule

module octaeightbitadd (
   input wire[31:0] a1,
   input wire[31:0] a2,
   input wire[31:0] a3,
   input wire[31:0] a4,
   input wire[31:0] a5,
   input wire[31:0] a6,
   input wire[31:0] a7,
   input wire[31:0] a8,
   input wire[31:0] b1,
   input wire[31:0] b2,
   input wire[31:0] b3,
   input wire[31:0] b4,
   input wire[31:0] b5,
   input wire[31:0] b6,
   input wire[31:0] b7,
   input wire[31:0] b8,
   output wire[31:0] sum,
   input clk,
);

reg [31:0] sum1;
reg [31:0] sum2;

 quadeightbitadd add1(
   .a1(a1),
   .a2(a2),
   .a3(a3),
   .a4(a4),
   .b1(a5),
   .b2(a6),
   .b3(a7),
   .b4(a8),
   .clk(clk),
   .sum(sum1),
);

 quadeightbitadd add2(
   .a1(b1),
   .a2(b2),
   .a3(b3),
   .a4(b4),
   .b1(b5),
   .b2(b6),
   .b3(b7),
   .b4(b8),
   .clk(clk),
   .sum(sum2),
);

 eightbitadd addTot(
   .a(sum1),
   .b(sum2),
   .c_in(1'b0),
   .clk(clk),
   .sum(sum),
);
endmodule

module hexaeightbitadd (
   input wire [31:0] a1,
   input wire [31:0] a2,
   input wire [31:0] a3,
   input wire [31:0] a4,
   input wire [31:0] a5,
   input wire [31:0] a6,
   input wire [31:0] a7,
   input wire [31:0] a8,
   input wire [31:0] a9,
   input wire [31:0] a10,
   input wire [31:0] a11,
   input wire [31:0] a12,
   input wire [31:0] a13,
   input wire [31:0] a14,
   input wire [31:0] a15,
   input wire [31:0] a16,
   input wire [31:0] b1,
   input wire [31:0] b2,
   input wire [31:0] b3,
   input wire [31:0] b4,
   input wire [31:0] b5,
   input wire [31:0] b6,
   input wire [31:0] b7,
   input wire [31:0] b8,
   input wire [31:0] b9,
   input wire [31:0] b10,
   input wire [31:0] b11,
   input wire [31:0] b12,
   input wire [31:0] b13,
   input wire [31:0] b14,
   input wire [31:0] b15,
   input wire [31:0] b16,
   output wire[31:0] sum,
   input clk,
);

reg [31:0] sum1;
reg [31:0] sum2;

 octaeightbitadd add1(
   .a1(a1),
   .a2(a2),
   .a3(a3),
   .a4(a4),
   .a5(a5),
   .a6(a6),
   .a7(a7),
   .a8(a8),
   .b1(a9),
   .b2(a10),
   .b3(a11),
   .b4(a12),
   .b5(a13),
   .b6(a14),
   .b7(a15),
   .b8(a16),
   .clk(clk),
   .sum(sum1),
);

 octaeightbitadd add2(
   .a1(b1),
   .a2(b2),
   .a3(b3),
   .a4(b4),
   .a5(b5),
   .a6(b6),
   .a7(b7),
   .a8(b8),
   .b1(b9),
   .b2(b10),
   .b3(b11),
   .b4(b12),
   .b5(b13),
   .b6(b14),
   .b7(b15),
   .b8(b16),
   .clk(clk),
   .sum(sum2),
);

 eightbitadd addTot(
   .a(sum1),
   .b(sum2),
   .c_in(1'b0),
   .clk(clk),
   .sum(sum),
);
endmodule


module activeTest(
   input inw,
   output outw,
);

// Initialize 48MHz clock
wire                                    CLK        ;
wire                                    CLK_RST    ;
reg         [31:0]                      counter    ;
reg         [31:0]                      sum        ;

reg outw;

qlal4s3b_cell_macro u_qlal4s3b_cell_macro (
    // FB Clocks
    .Sys_Clk0                  ( CLK                       ), // output
    .Sys_Clk0_Rst              ( CLK_RST                   ), // output
);

// Initialize Normal program
reg [31:0] v1;
reg [31:0] v2;
reg [31:0] v3;
reg [31:0] v4;
reg [31:0] v5;
reg [31:0] v6;
reg [31:0] v7;
reg [31:0] v8;
reg [31:0] v9;
reg [31:0] v10;
reg [31:0] v11;
reg [31:0] v12;
reg [31:0] v13;
reg [31:0] v14;
reg [31:0] v15;
reg [31:0] v16;
reg [31:0] v17;
reg [31:0] v18;
reg [31:0] v19;
reg [31:0] v20;
reg [31:0] v21;
reg [31:0] v22;
reg [31:0] v23;
reg [31:0] v24;
reg [31:0] v25;
reg [31:0] v26;
reg [31:0] v27;
reg [31:0] v28;
reg [31:0] v29;
reg [31:0] v30;
reg [31:0] v31;
reg [31:0] v32;

initial begin
   // Initialize values
   v1 <= 1;
   v2 <= 2;
   v3 <= 3;
   v4 <= 4;
   v5 <= 5;
   v6 <= 6;
   v7 <= 7;
   v8 <= 8;
   v9 <= 9;
   v10 <= 10;
   v11 <= 11;
   v12 <= 12;
   v13 <= 13;
   v14 <= 14;
   v15 <= 15;
   v16 <= 16;
   v17 <= 17;
   v18 <= 18;
   v19 <= 19;
   v20 <= 20;
   v21 <= 21;
   v22 <= 22;
   v23 <= 23;
   v24 <= 24;
   v25 <= 25;
   v26 <= 26;
   v27 <= 27;
   v28 <= 28;
   v29 <= 29;
   v30 <= 30;
   v31 <= 31;
   v32 <= 32;
   // Initialize counter
   counter <= 0;
end

hexaeightbitadd add1 (
   .a1(v1),
   .a2(v2),
   .a3(v3),
   .a4(v4),
   .a5(v5),
   .a6(v6),
   .a7(v7),
   .a8(v8),
   .a9(v9),
   .a10(v10),
   .a11(v11),
   .a12(v12),
   .a13(v13),
   .a14(v14),
   .a15(v15),
   .a16(v16),
   .b1(v17),
   .b2(v18),
   .b3(v19),
   .b4(v20),
   .b5(v21),
   .b6(v22),
   .b7(v23),
   .b8(v24),
   .b9(v25),
   .b10(v26),
   .b11(v27),
   .b12(v28),
   .b13(v29),
   .b14(v30),
   .b15(v31),
   .b16(v32),
   .sum(sum),
   .clk(CLK)
);

always @(posedge CLK) begin
   if (counter < 10000000) begin // Approx 1x every second
      counter <= counter + 1;
   end
   else begin
      if (inw) begin 
         v1 <= 1;
      end
      else begin
         v1 <= 30;
      end
      counter <= 0;
      if (sum == 528) begin // Check if correct value is computed
         outw <= 1;
      end
      else begin
         outw <= 0;
      end
   end
end
endmodule

module MODULE_top(
   io_pad
);

// GPIO
inout    wire     [31:0]      io_pad      ;

(*keep=1*)activeTest test (
   .inw(io_pad[6]),
   .outw(io_pad[21])
);

wire [1099:0] out;

reg en;
initial begin
   en <= 1;
end

lut_2_ro ro1(
   .en(en),
   .out(out[0]),
);

lut_2_ro ro2(
   .en(en),
   .out(out[1]),
);

lut_2_ro ro3(
   .en(en),
   .out(out[2]),
);

lut_2_ro ro4(
   .en(en),
   .out(out[3]),
);

lut_2_ro ro5(
   .en(en),
   .out(out[4]),
);

lut_2_ro ro6(
   .en(en),
   .out(out[5]),
);

lut_2_ro ro7(
   .en(en),
   .out(out[6]),
);

lut_2_ro ro8(
   .en(en),
   .out(out[7]),
);

lut_2_ro ro9(
   .en(en),
   .out(out[8]),
);

lut_2_ro ro10(
   .en(en),
   .out(out[9]),
);

lut_2_ro ro11(
   .en(en),
   .out(out[10]),
);

lut_2_ro ro12(
   .en(en),
   .out(out[11]),
);

lut_2_ro ro13(
   .en(en),
   .out(out[12]),
);

lut_2_ro ro14(
   .en(en),
   .out(out[13]),
);

lut_2_ro ro15(
   .en(en),
   .out(out[14]),
);

lut_2_ro ro16(
   .en(en),
   .out(out[15]),
);

lut_2_ro ro17(
   .en(en),
   .out(out[16]),
);

lut_2_ro ro18(
   .en(en),
   .out(out[17]),
);

lut_2_ro ro19(
   .en(en),
   .out(out[18]),
);

lut_2_ro ro20(
   .en(en),
   .out(out[19]),
);

lut_2_ro ro21(
   .en(en),
   .out(out[20]),
);

lut_2_ro ro22(
   .en(en),
   .out(out[21]),
);

lut_2_ro ro23(
   .en(en),
   .out(out[22]),
);

lut_2_ro ro24(
   .en(en),
   .out(out[23]),
);

lut_2_ro ro25(
   .en(en),
   .out(out[24]),
);

lut_2_ro ro26(
   .en(en),
   .out(out[25]),
);

lut_2_ro ro27(
   .en(en),
   .out(out[26]),
);

lut_2_ro ro28(
   .en(en),
   .out(out[27]),
);

lut_2_ro ro29(
   .en(en),
   .out(out[28]),
);

lut_2_ro ro30(
   .en(en),
   .out(out[29]),
);

lut_2_ro ro31(
   .en(en),
   .out(out[30]),
);

lut_2_ro ro32(
   .en(en),
   .out(out[31]),
);

lut_2_ro ro33(
   .en(en),
   .out(out[32]),
);

lut_2_ro ro34(
   .en(en),
   .out(out[33]),
);

lut_2_ro ro35(
   .en(en),
   .out(out[34]),
);

lut_2_ro ro36(
   .en(en),
   .out(out[35]),
);

lut_2_ro ro37(
   .en(en),
   .out(out[36]),
);

lut_2_ro ro38(
   .en(en),
   .out(out[37]),
);

lut_2_ro ro39(
   .en(en),
   .out(out[38]),
);

lut_2_ro ro40(
   .en(en),
   .out(out[39]),
);

lut_2_ro ro41(
   .en(en),
   .out(out[40]),
);

lut_2_ro ro42(
   .en(en),
   .out(out[41]),
);

lut_2_ro ro43(
   .en(en),
   .out(out[42]),
);

lut_2_ro ro44(
   .en(en),
   .out(out[43]),
);

lut_2_ro ro45(
   .en(en),
   .out(out[44]),
);

lut_2_ro ro46(
   .en(en),
   .out(out[45]),
);

lut_2_ro ro47(
   .en(en),
   .out(out[46]),
);

lut_2_ro ro48(
   .en(en),
   .out(out[47]),
);

lut_2_ro ro49(
   .en(en),
   .out(out[48]),
);

lut_2_ro ro50(
   .en(en),
   .out(out[49]),
);

lut_2_ro ro51(
   .en(en),
   .out(out[50]),
);

lut_2_ro ro52(
   .en(en),
   .out(out[51]),
);

lut_2_ro ro53(
   .en(en),
   .out(out[52]),
);

lut_2_ro ro54(
   .en(en),
   .out(out[53]),
);

lut_2_ro ro55(
   .en(en),
   .out(out[54]),
);

lut_2_ro ro56(
   .en(en),
   .out(out[55]),
);

lut_2_ro ro57(
   .en(en),
   .out(out[56]),
);

lut_2_ro ro58(
   .en(en),
   .out(out[57]),
);

lut_2_ro ro59(
   .en(en),
   .out(out[58]),
);

lut_2_ro ro60(
   .en(en),
   .out(out[59]),
);

lut_2_ro ro61(
   .en(en),
   .out(out[60]),
);

lut_2_ro ro62(
   .en(en),
   .out(out[61]),
);

lut_2_ro ro63(
   .en(en),
   .out(out[62]),
);

lut_2_ro ro64(
   .en(en),
   .out(out[63]),
);

lut_2_ro ro65(
   .en(en),
   .out(out[64]),
);

lut_2_ro ro66(
   .en(en),
   .out(out[65]),
);

lut_2_ro ro67(
   .en(en),
   .out(out[66]),
);

lut_2_ro ro68(
   .en(en),
   .out(out[67]),
);

lut_2_ro ro69(
   .en(en),
   .out(out[68]),
);

lut_2_ro ro70(
   .en(en),
   .out(out[69]),
);

lut_2_ro ro71(
   .en(en),
   .out(out[70]),
);

lut_2_ro ro72(
   .en(en),
   .out(out[71]),
);

lut_2_ro ro73(
   .en(en),
   .out(out[72]),
);

lut_2_ro ro74(
   .en(en),
   .out(out[73]),
);

lut_2_ro ro75(
   .en(en),
   .out(out[74]),
);

lut_2_ro ro76(
   .en(en),
   .out(out[75]),
);

lut_2_ro ro77(
   .en(en),
   .out(out[76]),
);

lut_2_ro ro78(
   .en(en),
   .out(out[77]),
);

lut_2_ro ro79(
   .en(en),
   .out(out[78]),
);

lut_2_ro ro80(
   .en(en),
   .out(out[79]),
);

lut_2_ro ro81(
   .en(en),
   .out(out[80]),
);

lut_2_ro ro82(
   .en(en),
   .out(out[81]),
);

lut_2_ro ro83(
   .en(en),
   .out(out[82]),
);

lut_2_ro ro84(
   .en(en),
   .out(out[83]),
);

lut_2_ro ro85(
   .en(en),
   .out(out[84]),
);

lut_2_ro ro86(
   .en(en),
   .out(out[85]),
);

lut_2_ro ro87(
   .en(en),
   .out(out[86]),
);

lut_2_ro ro88(
   .en(en),
   .out(out[87]),
);

lut_2_ro ro89(
   .en(en),
   .out(out[88]),
);

lut_2_ro ro90(
   .en(en),
   .out(out[89]),
);

lut_2_ro ro91(
   .en(en),
   .out(out[90]),
);

lut_2_ro ro92(
   .en(en),
   .out(out[91]),
);

lut_2_ro ro93(
   .en(en),
   .out(out[92]),
);

lut_2_ro ro94(
   .en(en),
   .out(out[93]),
);

lut_2_ro ro95(
   .en(en),
   .out(out[94]),
);

lut_2_ro ro96(
   .en(en),
   .out(out[95]),
);

lut_2_ro ro97(
   .en(en),
   .out(out[96]),
);

lut_2_ro ro98(
   .en(en),
   .out(out[97]),
);

lut_2_ro ro99(
   .en(en),
   .out(out[98]),
);

lut_2_ro ro100(
   .en(en),
   .out(out[99]),
);

lut_2_ro ro101(
   .en(en),
   .out(out[100]),
);

lut_2_ro ro102(
   .en(en),
   .out(out[101]),
);

lut_2_ro ro103(
   .en(en),
   .out(out[102]),
);

lut_2_ro ro104(
   .en(en),
   .out(out[103]),
);

lut_2_ro ro105(
   .en(en),
   .out(out[104]),
);

lut_2_ro ro106(
   .en(en),
   .out(out[105]),
);

lut_2_ro ro107(
   .en(en),
   .out(out[106]),
);

lut_2_ro ro108(
   .en(en),
   .out(out[107]),
);

lut_2_ro ro109(
   .en(en),
   .out(out[108]),
);

lut_2_ro ro110(
   .en(en),
   .out(out[109]),
);

lut_2_ro ro111(
   .en(en),
   .out(out[110]),
);

lut_2_ro ro112(
   .en(en),
   .out(out[111]),
);

lut_2_ro ro113(
   .en(en),
   .out(out[112]),
);

lut_2_ro ro114(
   .en(en),
   .out(out[113]),
);

lut_2_ro ro115(
   .en(en),
   .out(out[114]),
);

lut_2_ro ro116(
   .en(en),
   .out(out[115]),
);

lut_2_ro ro117(
   .en(en),
   .out(out[116]),
);

lut_2_ro ro118(
   .en(en),
   .out(out[117]),
);

lut_2_ro ro119(
   .en(en),
   .out(out[118]),
);

lut_2_ro ro120(
   .en(en),
   .out(out[119]),
);

lut_2_ro ro121(
   .en(en),
   .out(out[120]),
);

lut_2_ro ro122(
   .en(en),
   .out(out[121]),
);

lut_2_ro ro123(
   .en(en),
   .out(out[122]),
);

lut_2_ro ro124(
   .en(en),
   .out(out[123]),
);

lut_2_ro ro125(
   .en(en),
   .out(out[124]),
);

lut_2_ro ro126(
   .en(en),
   .out(out[125]),
);

lut_2_ro ro127(
   .en(en),
   .out(out[126]),
);

lut_2_ro ro128(
   .en(en),
   .out(out[127]),
);

lut_2_ro ro129(
   .en(en),
   .out(out[128]),
);

lut_2_ro ro130(
   .en(en),
   .out(out[129]),
);

lut_2_ro ro131(
   .en(en),
   .out(out[130]),
);

lut_2_ro ro132(
   .en(en),
   .out(out[131]),
);

lut_2_ro ro133(
   .en(en),
   .out(out[132]),
);

lut_2_ro ro134(
   .en(en),
   .out(out[133]),
);

lut_2_ro ro135(
   .en(en),
   .out(out[134]),
);

lut_2_ro ro136(
   .en(en),
   .out(out[135]),
);

lut_2_ro ro137(
   .en(en),
   .out(out[136]),
);

lut_2_ro ro138(
   .en(en),
   .out(out[137]),
);

lut_2_ro ro139(
   .en(en),
   .out(out[138]),
);

lut_2_ro ro140(
   .en(en),
   .out(out[139]),
);

lut_2_ro ro141(
   .en(en),
   .out(out[140]),
);

lut_2_ro ro142(
   .en(en),
   .out(out[141]),
);

lut_2_ro ro143(
   .en(en),
   .out(out[142]),
);

lut_2_ro ro144(
   .en(en),
   .out(out[143]),
);

lut_2_ro ro145(
   .en(en),
   .out(out[144]),
);

lut_2_ro ro146(
   .en(en),
   .out(out[145]),
);

lut_2_ro ro147(
   .en(en),
   .out(out[146]),
);

lut_2_ro ro148(
   .en(en),
   .out(out[147]),
);

lut_2_ro ro149(
   .en(en),
   .out(out[148]),
);

lut_2_ro ro150(
   .en(en),
   .out(out[149]),
);

lut_2_ro ro151(
   .en(en),
   .out(out[150]),
);

lut_2_ro ro152(
   .en(en),
   .out(out[151]),
);

lut_2_ro ro153(
   .en(en),
   .out(out[152]),
);

lut_2_ro ro154(
   .en(en),
   .out(out[153]),
);

lut_2_ro ro155(
   .en(en),
   .out(out[154]),
);

lut_2_ro ro156(
   .en(en),
   .out(out[155]),
);

lut_2_ro ro157(
   .en(en),
   .out(out[156]),
);

lut_2_ro ro158(
   .en(en),
   .out(out[157]),
);

lut_2_ro ro159(
   .en(en),
   .out(out[158]),
);

lut_2_ro ro160(
   .en(en),
   .out(out[159]),
);

lut_2_ro ro161(
   .en(en),
   .out(out[160]),
);

lut_2_ro ro162(
   .en(en),
   .out(out[161]),
);

lut_2_ro ro163(
   .en(en),
   .out(out[162]),
);

lut_2_ro ro164(
   .en(en),
   .out(out[163]),
);

lut_2_ro ro165(
   .en(en),
   .out(out[164]),
);

lut_2_ro ro166(
   .en(en),
   .out(out[165]),
);

lut_2_ro ro167(
   .en(en),
   .out(out[166]),
);

lut_2_ro ro168(
   .en(en),
   .out(out[167]),
);

lut_2_ro ro169(
   .en(en),
   .out(out[168]),
);

lut_2_ro ro170(
   .en(en),
   .out(out[169]),
);

lut_2_ro ro171(
   .en(en),
   .out(out[170]),
);

lut_2_ro ro172(
   .en(en),
   .out(out[171]),
);

lut_2_ro ro173(
   .en(en),
   .out(out[172]),
);

lut_2_ro ro174(
   .en(en),
   .out(out[173]),
);

lut_2_ro ro175(
   .en(en),
   .out(out[174]),
);

lut_2_ro ro176(
   .en(en),
   .out(out[175]),
);

lut_2_ro ro177(
   .en(en),
   .out(out[176]),
);

lut_2_ro ro178(
   .en(en),
   .out(out[177]),
);

lut_2_ro ro179(
   .en(en),
   .out(out[178]),
);

lut_2_ro ro180(
   .en(en),
   .out(out[179]),
);

lut_2_ro ro181(
   .en(en),
   .out(out[180]),
);

lut_2_ro ro182(
   .en(en),
   .out(out[181]),
);

lut_2_ro ro183(
   .en(en),
   .out(out[182]),
);

lut_2_ro ro184(
   .en(en),
   .out(out[183]),
);

lut_2_ro ro185(
   .en(en),
   .out(out[184]),
);

lut_2_ro ro186(
   .en(en),
   .out(out[185]),
);

lut_2_ro ro187(
   .en(en),
   .out(out[186]),
);

lut_2_ro ro188(
   .en(en),
   .out(out[187]),
);

lut_2_ro ro189(
   .en(en),
   .out(out[188]),
);

lut_2_ro ro190(
   .en(en),
   .out(out[189]),
);

lut_2_ro ro191(
   .en(en),
   .out(out[190]),
);

lut_2_ro ro192(
   .en(en),
   .out(out[191]),
);

lut_2_ro ro193(
   .en(en),
   .out(out[192]),
);

lut_2_ro ro194(
   .en(en),
   .out(out[193]),
);

lut_2_ro ro195(
   .en(en),
   .out(out[194]),
);

lut_2_ro ro196(
   .en(en),
   .out(out[195]),
);

lut_2_ro ro197(
   .en(en),
   .out(out[196]),
);

lut_2_ro ro198(
   .en(en),
   .out(out[197]),
);

lut_2_ro ro199(
   .en(en),
   .out(out[198]),
);

lut_2_ro ro200(
   .en(en),
   .out(out[199]),
);

lut_2_ro ro201(
   .en(en),
   .out(out[200]),
);

lut_2_ro ro202(
   .en(en),
   .out(out[201]),
);

lut_2_ro ro203(
   .en(en),
   .out(out[202]),
);

lut_2_ro ro204(
   .en(en),
   .out(out[203]),
);

lut_2_ro ro205(
   .en(en),
   .out(out[204]),
);

lut_2_ro ro206(
   .en(en),
   .out(out[205]),
);

lut_2_ro ro207(
   .en(en),
   .out(out[206]),
);

lut_2_ro ro208(
   .en(en),
   .out(out[207]),
);

lut_2_ro ro209(
   .en(en),
   .out(out[208]),
);

lut_2_ro ro210(
   .en(en),
   .out(out[209]),
);

lut_2_ro ro211(
   .en(en),
   .out(out[210]),
);

lut_2_ro ro212(
   .en(en),
   .out(out[211]),
);

lut_2_ro ro213(
   .en(en),
   .out(out[212]),
);

lut_2_ro ro214(
   .en(en),
   .out(out[213]),
);

lut_2_ro ro215(
   .en(en),
   .out(out[214]),
);

lut_2_ro ro216(
   .en(en),
   .out(out[215]),
);

lut_2_ro ro217(
   .en(en),
   .out(out[216]),
);

lut_2_ro ro218(
   .en(en),
   .out(out[217]),
);

lut_2_ro ro219(
   .en(en),
   .out(out[218]),
);

lut_2_ro ro220(
   .en(en),
   .out(out[219]),
);

lut_2_ro ro221(
   .en(en),
   .out(out[220]),
);

lut_2_ro ro222(
   .en(en),
   .out(out[221]),
);

lut_2_ro ro223(
   .en(en),
   .out(out[222]),
);

lut_2_ro ro224(
   .en(en),
   .out(out[223]),
);

lut_2_ro ro225(
   .en(en),
   .out(out[224]),
);

lut_2_ro ro226(
   .en(en),
   .out(out[225]),
);

lut_2_ro ro227(
   .en(en),
   .out(out[226]),
);

lut_2_ro ro228(
   .en(en),
   .out(out[227]),
);

lut_2_ro ro229(
   .en(en),
   .out(out[228]),
);

lut_2_ro ro230(
   .en(en),
   .out(out[229]),
);

lut_2_ro ro231(
   .en(en),
   .out(out[230]),
);

lut_2_ro ro232(
   .en(en),
   .out(out[231]),
);

lut_2_ro ro233(
   .en(en),
   .out(out[232]),
);

lut_2_ro ro234(
   .en(en),
   .out(out[233]),
);

lut_2_ro ro235(
   .en(en),
   .out(out[234]),
);

lut_2_ro ro236(
   .en(en),
   .out(out[235]),
);

lut_2_ro ro237(
   .en(en),
   .out(out[236]),
);

lut_2_ro ro238(
   .en(en),
   .out(out[237]),
);

lut_2_ro ro239(
   .en(en),
   .out(out[238]),
);

lut_2_ro ro240(
   .en(en),
   .out(out[239]),
);

lut_2_ro ro241(
   .en(en),
   .out(out[240]),
);

lut_2_ro ro242(
   .en(en),
   .out(out[241]),
);

lut_2_ro ro243(
   .en(en),
   .out(out[242]),
);

lut_2_ro ro244(
   .en(en),
   .out(out[243]),
);

lut_2_ro ro245(
   .en(en),
   .out(out[244]),
);

lut_2_ro ro246(
   .en(en),
   .out(out[245]),
);

lut_2_ro ro247(
   .en(en),
   .out(out[246]),
);

lut_2_ro ro248(
   .en(en),
   .out(out[247]),
);

lut_2_ro ro249(
   .en(en),
   .out(out[248]),
);

lut_2_ro ro250(
   .en(en),
   .out(out[249]),
);

lut_2_ro ro251(
   .en(en),
   .out(out[250]),
);

lut_2_ro ro252(
   .en(en),
   .out(out[251]),
);

lut_2_ro ro253(
   .en(en),
   .out(out[252]),
);

lut_2_ro ro254(
   .en(en),
   .out(out[253]),
);

lut_2_ro ro255(
   .en(en),
   .out(out[254]),
);

lut_2_ro ro256(
   .en(en),
   .out(out[255]),
);

lut_2_ro ro257(
   .en(en),
   .out(out[256]),
);

lut_2_ro ro258(
   .en(en),
   .out(out[257]),
);

lut_2_ro ro259(
   .en(en),
   .out(out[258]),
);

lut_2_ro ro260(
   .en(en),
   .out(out[259]),
);

lut_2_ro ro261(
   .en(en),
   .out(out[260]),
);

lut_2_ro ro262(
   .en(en),
   .out(out[261]),
);

lut_2_ro ro263(
   .en(en),
   .out(out[262]),
);

lut_2_ro ro264(
   .en(en),
   .out(out[263]),
);

lut_2_ro ro265(
   .en(en),
   .out(out[264]),
);

lut_2_ro ro266(
   .en(en),
   .out(out[265]),
);

lut_2_ro ro267(
   .en(en),
   .out(out[266]),
);

lut_2_ro ro268(
   .en(en),
   .out(out[267]),
);

lut_2_ro ro269(
   .en(en),
   .out(out[268]),
);

lut_2_ro ro270(
   .en(en),
   .out(out[269]),
);

lut_2_ro ro271(
   .en(en),
   .out(out[270]),
);

lut_2_ro ro272(
   .en(en),
   .out(out[271]),
);

lut_2_ro ro273(
   .en(en),
   .out(out[272]),
);

lut_2_ro ro274(
   .en(en),
   .out(out[273]),
);

lut_2_ro ro275(
   .en(en),
   .out(out[274]),
);

lut_2_ro ro276(
   .en(en),
   .out(out[275]),
);

lut_2_ro ro277(
   .en(en),
   .out(out[276]),
);

lut_2_ro ro278(
   .en(en),
   .out(out[277]),
);

lut_2_ro ro279(
   .en(en),
   .out(out[278]),
);

lut_2_ro ro280(
   .en(en),
   .out(out[279]),
);

lut_2_ro ro281(
   .en(en),
   .out(out[280]),
);

lut_2_ro ro282(
   .en(en),
   .out(out[281]),
);

lut_2_ro ro283(
   .en(en),
   .out(out[282]),
);

lut_2_ro ro284(
   .en(en),
   .out(out[283]),
);

lut_2_ro ro285(
   .en(en),
   .out(out[284]),
);

lut_2_ro ro286(
   .en(en),
   .out(out[285]),
);

lut_2_ro ro287(
   .en(en),
   .out(out[286]),
);

lut_2_ro ro288(
   .en(en),
   .out(out[287]),
);

lut_2_ro ro289(
   .en(en),
   .out(out[288]),
);

lut_2_ro ro290(
   .en(en),
   .out(out[289]),
);

lut_2_ro ro291(
   .en(en),
   .out(out[290]),
);

lut_2_ro ro292(
   .en(en),
   .out(out[291]),
);

lut_2_ro ro293(
   .en(en),
   .out(out[292]),
);

lut_2_ro ro294(
   .en(en),
   .out(out[293]),
);

lut_2_ro ro295(
   .en(en),
   .out(out[294]),
);

lut_2_ro ro296(
   .en(en),
   .out(out[295]),
);

lut_2_ro ro297(
   .en(en),
   .out(out[296]),
);

lut_2_ro ro298(
   .en(en),
   .out(out[297]),
);

lut_2_ro ro299(
   .en(en),
   .out(out[298]),
);

lut_2_ro ro300(
   .en(en),
   .out(out[299]),
);

lut_2_ro ro301(
   .en(en),
   .out(out[300]),
);

lut_2_ro ro302(
   .en(en),
   .out(out[301]),
);

lut_2_ro ro303(
   .en(en),
   .out(out[302]),
);

lut_2_ro ro304(
   .en(en),
   .out(out[303]),
);

lut_2_ro ro305(
   .en(en),
   .out(out[304]),
);

lut_2_ro ro306(
   .en(en),
   .out(out[305]),
);

lut_2_ro ro307(
   .en(en),
   .out(out[306]),
);

lut_2_ro ro308(
   .en(en),
   .out(out[307]),
);

lut_2_ro ro309(
   .en(en),
   .out(out[308]),
);

lut_2_ro ro310(
   .en(en),
   .out(out[309]),
);

lut_2_ro ro311(
   .en(en),
   .out(out[310]),
);

lut_2_ro ro312(
   .en(en),
   .out(out[311]),
);

lut_2_ro ro313(
   .en(en),
   .out(out[312]),
);

lut_2_ro ro314(
   .en(en),
   .out(out[313]),
);

lut_2_ro ro315(
   .en(en),
   .out(out[314]),
);

lut_2_ro ro316(
   .en(en),
   .out(out[315]),
);

lut_2_ro ro317(
   .en(en),
   .out(out[316]),
);

lut_2_ro ro318(
   .en(en),
   .out(out[317]),
);

lut_2_ro ro319(
   .en(en),
   .out(out[318]),
);

lut_2_ro ro320(
   .en(en),
   .out(out[319]),
);

lut_2_ro ro321(
   .en(en),
   .out(out[320]),
);

lut_2_ro ro322(
   .en(en),
   .out(out[321]),
);

lut_2_ro ro323(
   .en(en),
   .out(out[322]),
);

lut_2_ro ro324(
   .en(en),
   .out(out[323]),
);

lut_2_ro ro325(
   .en(en),
   .out(out[324]),
);

lut_2_ro ro326(
   .en(en),
   .out(out[325]),
);

lut_2_ro ro327(
   .en(en),
   .out(out[326]),
);

lut_2_ro ro328(
   .en(en),
   .out(out[327]),
);

lut_2_ro ro329(
   .en(en),
   .out(out[328]),
);

lut_2_ro ro330(
   .en(en),
   .out(out[329]),
);

lut_2_ro ro331(
   .en(en),
   .out(out[330]),
);

lut_2_ro ro332(
   .en(en),
   .out(out[331]),
);

lut_2_ro ro333(
   .en(en),
   .out(out[332]),
);

lut_2_ro ro334(
   .en(en),
   .out(out[333]),
);

lut_2_ro ro335(
   .en(en),
   .out(out[334]),
);

lut_2_ro ro336(
   .en(en),
   .out(out[335]),
);

lut_2_ro ro337(
   .en(en),
   .out(out[336]),
);

lut_2_ro ro338(
   .en(en),
   .out(out[337]),
);

lut_2_ro ro339(
   .en(en),
   .out(out[338]),
);

lut_2_ro ro340(
   .en(en),
   .out(out[339]),
);

lut_2_ro ro341(
   .en(en),
   .out(out[340]),
);

lut_2_ro ro342(
   .en(en),
   .out(out[341]),
);

lut_2_ro ro343(
   .en(en),
   .out(out[342]),
);

lut_2_ro ro344(
   .en(en),
   .out(out[343]),
);

lut_2_ro ro345(
   .en(en),
   .out(out[344]),
);

lut_2_ro ro346(
   .en(en),
   .out(out[345]),
);

lut_2_ro ro347(
   .en(en),
   .out(out[346]),
);

lut_2_ro ro348(
   .en(en),
   .out(out[347]),
);

lut_2_ro ro349(
   .en(en),
   .out(out[348]),
);

lut_2_ro ro350(
   .en(en),
   .out(out[349]),
);

lut_2_ro ro351(
   .en(en),
   .out(out[350]),
);

lut_2_ro ro352(
   .en(en),
   .out(out[351]),
);

lut_2_ro ro353(
   .en(en),
   .out(out[352]),
);

lut_2_ro ro354(
   .en(en),
   .out(out[353]),
);

lut_2_ro ro355(
   .en(en),
   .out(out[354]),
);

lut_2_ro ro356(
   .en(en),
   .out(out[355]),
);

lut_2_ro ro357(
   .en(en),
   .out(out[356]),
);

lut_2_ro ro358(
   .en(en),
   .out(out[357]),
);

lut_2_ro ro359(
   .en(en),
   .out(out[358]),
);

lut_2_ro ro360(
   .en(en),
   .out(out[359]),
);

lut_2_ro ro361(
   .en(en),
   .out(out[360]),
);

lut_2_ro ro362(
   .en(en),
   .out(out[361]),
);

lut_2_ro ro363(
   .en(en),
   .out(out[362]),
);

lut_2_ro ro364(
   .en(en),
   .out(out[363]),
);

lut_2_ro ro365(
   .en(en),
   .out(out[364]),
);

lut_2_ro ro366(
   .en(en),
   .out(out[365]),
);

lut_2_ro ro367(
   .en(en),
   .out(out[366]),
);

lut_2_ro ro368(
   .en(en),
   .out(out[367]),
);

lut_2_ro ro369(
   .en(en),
   .out(out[368]),
);

lut_2_ro ro370(
   .en(en),
   .out(out[369]),
);

lut_2_ro ro371(
   .en(en),
   .out(out[370]),
);

lut_2_ro ro372(
   .en(en),
   .out(out[371]),
);

lut_2_ro ro373(
   .en(en),
   .out(out[372]),
);

lut_2_ro ro374(
   .en(en),
   .out(out[373]),
);

lut_2_ro ro375(
   .en(en),
   .out(out[374]),
);

lut_2_ro ro376(
   .en(en),
   .out(out[375]),
);

lut_2_ro ro377(
   .en(en),
   .out(out[376]),
);

lut_2_ro ro378(
   .en(en),
   .out(out[377]),
);

lut_2_ro ro379(
   .en(en),
   .out(out[378]),
);

lut_2_ro ro380(
   .en(en),
   .out(out[379]),
);

lut_2_ro ro381(
   .en(en),
   .out(out[380]),
);

lut_2_ro ro382(
   .en(en),
   .out(out[381]),
);

lut_2_ro ro383(
   .en(en),
   .out(out[382]),
);

lut_2_ro ro384(
   .en(en),
   .out(out[383]),
);

lut_2_ro ro385(
   .en(en),
   .out(out[384]),
);

lut_2_ro ro386(
   .en(en),
   .out(out[385]),
);

lut_2_ro ro387(
   .en(en),
   .out(out[386]),
);

lut_2_ro ro388(
   .en(en),
   .out(out[387]),
);

lut_2_ro ro389(
   .en(en),
   .out(out[388]),
);

lut_2_ro ro390(
   .en(en),
   .out(out[389]),
);

lut_2_ro ro391(
   .en(en),
   .out(out[390]),
);

lut_2_ro ro392(
   .en(en),
   .out(out[391]),
);

lut_2_ro ro393(
   .en(en),
   .out(out[392]),
);

lut_2_ro ro394(
   .en(en),
   .out(out[393]),
);

lut_2_ro ro395(
   .en(en),
   .out(out[394]),
);

lut_2_ro ro396(
   .en(en),
   .out(out[395]),
);

lut_2_ro ro397(
   .en(en),
   .out(out[396]),
);

lut_2_ro ro398(
   .en(en),
   .out(out[397]),
);

lut_2_ro ro399(
   .en(en),
   .out(out[398]),
);

lut_2_ro ro400(
   .en(en),
   .out(out[399]),
);

lut_2_ro ro401(
   .en(en),
   .out(out[400]),
);

lut_2_ro ro402(
   .en(en),
   .out(out[401]),
);

lut_2_ro ro403(
   .en(en),
   .out(out[402]),
);

lut_2_ro ro404(
   .en(en),
   .out(out[403]),
);

lut_2_ro ro405(
   .en(en),
   .out(out[404]),
);

lut_2_ro ro406(
   .en(en),
   .out(out[405]),
);

lut_2_ro ro407(
   .en(en),
   .out(out[406]),
);

lut_2_ro ro408(
   .en(en),
   .out(out[407]),
);

lut_2_ro ro409(
   .en(en),
   .out(out[408]),
);

lut_2_ro ro410(
   .en(en),
   .out(out[409]),
);

lut_2_ro ro411(
   .en(en),
   .out(out[410]),
);

lut_2_ro ro412(
   .en(en),
   .out(out[411]),
);

lut_2_ro ro413(
   .en(en),
   .out(out[412]),
);

lut_2_ro ro414(
   .en(en),
   .out(out[413]),
);

lut_2_ro ro415(
   .en(en),
   .out(out[414]),
);

lut_2_ro ro416(
   .en(en),
   .out(out[415]),
);

lut_2_ro ro417(
   .en(en),
   .out(out[416]),
);

lut_2_ro ro418(
   .en(en),
   .out(out[417]),
);

lut_2_ro ro419(
   .en(en),
   .out(out[418]),
);

lut_2_ro ro420(
   .en(en),
   .out(out[419]),
);

lut_2_ro ro421(
   .en(en),
   .out(out[420]),
);

lut_2_ro ro422(
   .en(en),
   .out(out[421]),
);

lut_2_ro ro423(
   .en(en),
   .out(out[422]),
);

lut_2_ro ro424(
   .en(en),
   .out(out[423]),
);

lut_2_ro ro425(
   .en(en),
   .out(out[424]),
);

lut_2_ro ro426(
   .en(en),
   .out(out[425]),
);

lut_2_ro ro427(
   .en(en),
   .out(out[426]),
);

lut_2_ro ro428(
   .en(en),
   .out(out[427]),
);

lut_2_ro ro429(
   .en(en),
   .out(out[428]),
);

lut_2_ro ro430(
   .en(en),
   .out(out[429]),
);

lut_2_ro ro431(
   .en(en),
   .out(out[430]),
);

lut_2_ro ro432(
   .en(en),
   .out(out[431]),
);

lut_2_ro ro433(
   .en(en),
   .out(out[432]),
);

lut_2_ro ro434(
   .en(en),
   .out(out[433]),
);

lut_2_ro ro435(
   .en(en),
   .out(out[434]),
);

lut_2_ro ro436(
   .en(en),
   .out(out[435]),
);

lut_2_ro ro437(
   .en(en),
   .out(out[436]),
);

lut_2_ro ro438(
   .en(en),
   .out(out[437]),
);

lut_2_ro ro439(
   .en(en),
   .out(out[438]),
);

lut_2_ro ro440(
   .en(en),
   .out(out[439]),
);

lut_2_ro ro441(
   .en(en),
   .out(out[440]),
);

lut_2_ro ro442(
   .en(en),
   .out(out[441]),
);

lut_2_ro ro443(
   .en(en),
   .out(out[442]),
);

lut_2_ro ro444(
   .en(en),
   .out(out[443]),
);

lut_2_ro ro445(
   .en(en),
   .out(out[444]),
);

lut_2_ro ro446(
   .en(en),
   .out(out[445]),
);

lut_2_ro ro447(
   .en(en),
   .out(out[446]),
);

lut_2_ro ro448(
   .en(en),
   .out(out[447]),
);

lut_2_ro ro449(
   .en(en),
   .out(out[448]),
);

lut_2_ro ro450(
   .en(en),
   .out(out[449]),
);

lut_2_ro ro451(
   .en(en),
   .out(out[450]),
);

lut_2_ro ro452(
   .en(en),
   .out(out[451]),
);

lut_2_ro ro453(
   .en(en),
   .out(out[452]),
);

lut_2_ro ro454(
   .en(en),
   .out(out[453]),
);

lut_2_ro ro455(
   .en(en),
   .out(out[454]),
);

lut_2_ro ro456(
   .en(en),
   .out(out[455]),
);

lut_2_ro ro457(
   .en(en),
   .out(out[456]),
);

lut_2_ro ro458(
   .en(en),
   .out(out[457]),
);

lut_2_ro ro459(
   .en(en),
   .out(out[458]),
);

lut_2_ro ro460(
   .en(en),
   .out(out[459]),
);

lut_2_ro ro461(
   .en(en),
   .out(out[460]),
);

lut_2_ro ro462(
   .en(en),
   .out(out[461]),
);

lut_2_ro ro463(
   .en(en),
   .out(out[462]),
);

lut_2_ro ro464(
   .en(en),
   .out(out[463]),
);

lut_2_ro ro465(
   .en(en),
   .out(out[464]),
);

lut_2_ro ro466(
   .en(en),
   .out(out[465]),
);

lut_2_ro ro467(
   .en(en),
   .out(out[466]),
);

lut_2_ro ro468(
   .en(en),
   .out(out[467]),
);

lut_2_ro ro469(
   .en(en),
   .out(out[468]),
);

lut_2_ro ro470(
   .en(en),
   .out(out[469]),
);

lut_2_ro ro471(
   .en(en),
   .out(out[470]),
);

lut_2_ro ro472(
   .en(en),
   .out(out[471]),
);

lut_2_ro ro473(
   .en(en),
   .out(out[472]),
);

lut_2_ro ro474(
   .en(en),
   .out(out[473]),
);

lut_2_ro ro475(
   .en(en),
   .out(out[474]),
);

lut_2_ro ro476(
   .en(en),
   .out(out[475]),
);

lut_2_ro ro477(
   .en(en),
   .out(out[476]),
);

lut_2_ro ro478(
   .en(en),
   .out(out[477]),
);

lut_2_ro ro479(
   .en(en),
   .out(out[478]),
);

lut_2_ro ro480(
   .en(en),
   .out(out[479]),
);

lut_2_ro ro481(
   .en(en),
   .out(out[480]),
);

lut_2_ro ro482(
   .en(en),
   .out(out[481]),
);

lut_2_ro ro483(
   .en(en),
   .out(out[482]),
);

lut_2_ro ro484(
   .en(en),
   .out(out[483]),
);

lut_2_ro ro485(
   .en(en),
   .out(out[484]),
);

lut_2_ro ro486(
   .en(en),
   .out(out[485]),
);

lut_2_ro ro487(
   .en(en),
   .out(out[486]),
);

lut_2_ro ro488(
   .en(en),
   .out(out[487]),
);

lut_2_ro ro489(
   .en(en),
   .out(out[488]),
);

lut_2_ro ro490(
   .en(en),
   .out(out[489]),
);

lut_2_ro ro491(
   .en(en),
   .out(out[490]),
);

lut_2_ro ro492(
   .en(en),
   .out(out[491]),
);

lut_2_ro ro493(
   .en(en),
   .out(out[492]),
);

lut_2_ro ro494(
   .en(en),
   .out(out[493]),
);

lut_2_ro ro495(
   .en(en),
   .out(out[494]),
);

lut_2_ro ro496(
   .en(en),
   .out(out[495]),
);

lut_2_ro ro497(
   .en(en),
   .out(out[496]),
);

lut_2_ro ro498(
   .en(en),
   .out(out[497]),
);

lut_2_ro ro499(
   .en(en),
   .out(out[498]),
);

lut_2_ro ro500(
   .en(en),
   .out(out[499]),
);

lut_2_ro ro501(
   .en(en),
   .out(out[500]),
);

lut_2_ro ro502(
   .en(en),
   .out(out[501]),
);

lut_2_ro ro503(
   .en(en),
   .out(out[502]),
);

lut_2_ro ro504(
   .en(en),
   .out(out[503]),
);

lut_2_ro ro505(
   .en(en),
   .out(out[504]),
);

lut_2_ro ro506(
   .en(en),
   .out(out[505]),
);

lut_2_ro ro507(
   .en(en),
   .out(out[506]),
);

lut_2_ro ro508(
   .en(en),
   .out(out[507]),
);

lut_2_ro ro509(
   .en(en),
   .out(out[508]),
);

lut_2_ro ro510(
   .en(en),
   .out(out[509]),
);

lut_2_ro ro511(
   .en(en),
   .out(out[510]),
);

lut_2_ro ro512(
   .en(en),
   .out(out[511]),
);

lut_2_ro ro513(
   .en(en),
   .out(out[512]),
);

lut_2_ro ro514(
   .en(en),
   .out(out[513]),
);

lut_2_ro ro515(
   .en(en),
   .out(out[514]),
);

lut_2_ro ro516(
   .en(en),
   .out(out[515]),
);

lut_2_ro ro517(
   .en(en),
   .out(out[516]),
);

lut_2_ro ro518(
   .en(en),
   .out(out[517]),
);

lut_2_ro ro519(
   .en(en),
   .out(out[518]),
);

lut_2_ro ro520(
   .en(en),
   .out(out[519]),
);

lut_2_ro ro521(
   .en(en),
   .out(out[520]),
);

lut_2_ro ro522(
   .en(en),
   .out(out[521]),
);

lut_2_ro ro523(
   .en(en),
   .out(out[522]),
);

lut_2_ro ro524(
   .en(en),
   .out(out[523]),
);

lut_2_ro ro525(
   .en(en),
   .out(out[524]),
);

lut_2_ro ro526(
   .en(en),
   .out(out[525]),
);

lut_2_ro ro527(
   .en(en),
   .out(out[526]),
);

lut_2_ro ro528(
   .en(en),
   .out(out[527]),
);

lut_2_ro ro529(
   .en(en),
   .out(out[528]),
);

lut_2_ro ro530(
   .en(en),
   .out(out[529]),
);

lut_2_ro ro531(
   .en(en),
   .out(out[530]),
);

lut_2_ro ro532(
   .en(en),
   .out(out[531]),
);

lut_2_ro ro533(
   .en(en),
   .out(out[532]),
);

lut_2_ro ro534(
   .en(en),
   .out(out[533]),
);

lut_2_ro ro535(
   .en(en),
   .out(out[534]),
);

lut_2_ro ro536(
   .en(en),
   .out(out[535]),
);

lut_2_ro ro537(
   .en(en),
   .out(out[536]),
);

lut_2_ro ro538(
   .en(en),
   .out(out[537]),
);

lut_2_ro ro539(
   .en(en),
   .out(out[538]),
);

lut_2_ro ro540(
   .en(en),
   .out(out[539]),
);

lut_2_ro ro541(
   .en(en),
   .out(out[540]),
);

lut_2_ro ro542(
   .en(en),
   .out(out[541]),
);

lut_2_ro ro543(
   .en(en),
   .out(out[542]),
);

lut_2_ro ro544(
   .en(en),
   .out(out[543]),
);

lut_2_ro ro545(
   .en(en),
   .out(out[544]),
);

lut_2_ro ro546(
   .en(en),
   .out(out[545]),
);

lut_2_ro ro547(
   .en(en),
   .out(out[546]),
);

lut_2_ro ro548(
   .en(en),
   .out(out[547]),
);

lut_2_ro ro549(
   .en(en),
   .out(out[548]),
);

lut_2_ro ro550(
   .en(en),
   .out(out[549]),
);

lut_2_ro ro551(
   .en(en),
   .out(out[550]),
);

lut_2_ro ro552(
   .en(en),
   .out(out[551]),
);

lut_2_ro ro553(
   .en(en),
   .out(out[552]),
);

lut_2_ro ro554(
   .en(en),
   .out(out[553]),
);

lut_2_ro ro555(
   .en(en),
   .out(out[554]),
);

lut_2_ro ro556(
   .en(en),
   .out(out[555]),
);

lut_2_ro ro557(
   .en(en),
   .out(out[556]),
);

lut_2_ro ro558(
   .en(en),
   .out(out[557]),
);

lut_2_ro ro559(
   .en(en),
   .out(out[558]),
);

lut_2_ro ro560(
   .en(en),
   .out(out[559]),
);

lut_2_ro ro561(
   .en(en),
   .out(out[560]),
);

lut_2_ro ro562(
   .en(en),
   .out(out[561]),
);

lut_2_ro ro563(
   .en(en),
   .out(out[562]),
);

lut_2_ro ro564(
   .en(en),
   .out(out[563]),
);

lut_2_ro ro565(
   .en(en),
   .out(out[564]),
);

lut_2_ro ro566(
   .en(en),
   .out(out[565]),
);

lut_2_ro ro567(
   .en(en),
   .out(out[566]),
);

lut_2_ro ro568(
   .en(en),
   .out(out[567]),
);

lut_2_ro ro569(
   .en(en),
   .out(out[568]),
);

lut_2_ro ro570(
   .en(en),
   .out(out[569]),
);

lut_2_ro ro571(
   .en(en),
   .out(out[570]),
);

lut_2_ro ro572(
   .en(en),
   .out(out[571]),
);

lut_2_ro ro573(
   .en(en),
   .out(out[572]),
);

lut_2_ro ro574(
   .en(en),
   .out(out[573]),
);

lut_2_ro ro575(
   .en(en),
   .out(out[574]),
);

lut_2_ro ro576(
   .en(en),
   .out(out[575]),
);

lut_2_ro ro577(
   .en(en),
   .out(out[576]),
);

lut_2_ro ro578(
   .en(en),
   .out(out[577]),
);

lut_2_ro ro579(
   .en(en),
   .out(out[578]),
);

lut_2_ro ro580(
   .en(en),
   .out(out[579]),
);

lut_2_ro ro581(
   .en(en),
   .out(out[580]),
);

lut_2_ro ro582(
   .en(en),
   .out(out[581]),
);

lut_2_ro ro583(
   .en(en),
   .out(out[582]),
);

lut_2_ro ro584(
   .en(en),
   .out(out[583]),
);

lut_2_ro ro585(
   .en(en),
   .out(out[584]),
);

lut_2_ro ro586(
   .en(en),
   .out(out[585]),
);

lut_2_ro ro587(
   .en(en),
   .out(out[586]),
);

lut_2_ro ro588(
   .en(en),
   .out(out[587]),
);

lut_2_ro ro589(
   .en(en),
   .out(out[588]),
);

lut_2_ro ro590(
   .en(en),
   .out(out[589]),
);

lut_2_ro ro591(
   .en(en),
   .out(out[590]),
);

lut_2_ro ro592(
   .en(en),
   .out(out[591]),
);

lut_2_ro ro593(
   .en(en),
   .out(out[592]),
);

lut_2_ro ro594(
   .en(en),
   .out(out[593]),
);

lut_2_ro ro595(
   .en(en),
   .out(out[594]),
);

lut_2_ro ro596(
   .en(en),
   .out(out[595]),
);

lut_2_ro ro597(
   .en(en),
   .out(out[596]),
);

lut_2_ro ro598(
   .en(en),
   .out(out[597]),
);

lut_2_ro ro599(
   .en(en),
   .out(out[598]),
);

lut_2_ro ro600(
   .en(en),
   .out(out[599]),
);

lut_2_ro ro601(
   .en(en),
   .out(out[600]),
);

lut_2_ro ro602(
   .en(en),
   .out(out[601]),
);

lut_2_ro ro603(
   .en(en),
   .out(out[602]),
);

lut_2_ro ro604(
   .en(en),
   .out(out[603]),
);

lut_2_ro ro605(
   .en(en),
   .out(out[604]),
);

lut_2_ro ro606(
   .en(en),
   .out(out[605]),
);

lut_2_ro ro607(
   .en(en),
   .out(out[606]),
);

lut_2_ro ro608(
   .en(en),
   .out(out[607]),
);

lut_2_ro ro609(
   .en(en),
   .out(out[608]),
);

lut_2_ro ro610(
   .en(en),
   .out(out[609]),
);

lut_2_ro ro611(
   .en(en),
   .out(out[610]),
);

lut_2_ro ro612(
   .en(en),
   .out(out[611]),
);

lut_2_ro ro613(
   .en(en),
   .out(out[612]),
);

lut_2_ro ro614(
   .en(en),
   .out(out[613]),
);

lut_2_ro ro615(
   .en(en),
   .out(out[614]),
);

lut_2_ro ro616(
   .en(en),
   .out(out[615]),
);

lut_2_ro ro617(
   .en(en),
   .out(out[616]),
);

lut_2_ro ro618(
   .en(en),
   .out(out[617]),
);

lut_2_ro ro619(
   .en(en),
   .out(out[618]),
);

lut_2_ro ro620(
   .en(en),
   .out(out[619]),
);

lut_2_ro ro621(
   .en(en),
   .out(out[620]),
);

lut_2_ro ro622(
   .en(en),
   .out(out[621]),
);

lut_2_ro ro623(
   .en(en),
   .out(out[622]),
);

lut_2_ro ro624(
   .en(en),
   .out(out[623]),
);

lut_2_ro ro625(
   .en(en),
   .out(out[624]),
);

lut_2_ro ro626(
   .en(en),
   .out(out[625]),
);

lut_2_ro ro627(
   .en(en),
   .out(out[626]),
);

lut_2_ro ro628(
   .en(en),
   .out(out[627]),
);

lut_2_ro ro629(
   .en(en),
   .out(out[628]),
);

lut_2_ro ro630(
   .en(en),
   .out(out[629]),
);

lut_2_ro ro631(
   .en(en),
   .out(out[630]),
);

lut_2_ro ro632(
   .en(en),
   .out(out[631]),
);

lut_2_ro ro633(
   .en(en),
   .out(out[632]),
);

lut_2_ro ro634(
   .en(en),
   .out(out[633]),
);

lut_2_ro ro635(
   .en(en),
   .out(out[634]),
);

lut_2_ro ro636(
   .en(en),
   .out(out[635]),
);

lut_2_ro ro637(
   .en(en),
   .out(out[636]),
);

lut_2_ro ro638(
   .en(en),
   .out(out[637]),
);

lut_2_ro ro639(
   .en(en),
   .out(out[638]),
);

lut_2_ro ro640(
   .en(en),
   .out(out[639]),
);

lut_2_ro ro641(
   .en(en),
   .out(out[640]),
);

lut_2_ro ro642(
   .en(en),
   .out(out[641]),
);

lut_2_ro ro643(
   .en(en),
   .out(out[642]),
);

lut_2_ro ro644(
   .en(en),
   .out(out[643]),
);

lut_2_ro ro645(
   .en(en),
   .out(out[644]),
);

lut_2_ro ro646(
   .en(en),
   .out(out[645]),
);

lut_2_ro ro647(
   .en(en),
   .out(out[646]),
);

lut_2_ro ro648(
   .en(en),
   .out(out[647]),
);

lut_2_ro ro649(
   .en(en),
   .out(out[648]),
);

lut_2_ro ro650(
   .en(en),
   .out(out[649]),
);

lut_2_ro ro651(
   .en(en),
   .out(out[650]),
);

lut_2_ro ro652(
   .en(en),
   .out(out[651]),
);

lut_2_ro ro653(
   .en(en),
   .out(out[652]),
);

lut_2_ro ro654(
   .en(en),
   .out(out[653]),
);

lut_2_ro ro655(
   .en(en),
   .out(out[654]),
);

lut_2_ro ro656(
   .en(en),
   .out(out[655]),
);

lut_2_ro ro657(
   .en(en),
   .out(out[656]),
);

lut_2_ro ro658(
   .en(en),
   .out(out[657]),
);

lut_2_ro ro659(
   .en(en),
   .out(out[658]),
);

lut_2_ro ro660(
   .en(en),
   .out(out[659]),
);

lut_2_ro ro661(
   .en(en),
   .out(out[660]),
);

lut_2_ro ro662(
   .en(en),
   .out(out[661]),
);

lut_2_ro ro663(
   .en(en),
   .out(out[662]),
);

lut_2_ro ro664(
   .en(en),
   .out(out[663]),
);

lut_2_ro ro665(
   .en(en),
   .out(out[664]),
);

lut_2_ro ro666(
   .en(en),
   .out(out[665]),
);

lut_2_ro ro667(
   .en(en),
   .out(out[666]),
);

lut_2_ro ro668(
   .en(en),
   .out(out[667]),
);

lut_2_ro ro669(
   .en(en),
   .out(out[668]),
);

lut_2_ro ro670(
   .en(en),
   .out(out[669]),
);

lut_2_ro ro671(
   .en(en),
   .out(out[670]),
);

lut_2_ro ro672(
   .en(en),
   .out(out[671]),
);

lut_2_ro ro673(
   .en(en),
   .out(out[672]),
);

lut_2_ro ro674(
   .en(en),
   .out(out[673]),
);

lut_2_ro ro675(
   .en(en),
   .out(out[674]),
);

lut_2_ro ro676(
   .en(en),
   .out(out[675]),
);

lut_2_ro ro677(
   .en(en),
   .out(out[676]),
);

lut_2_ro ro678(
   .en(en),
   .out(out[677]),
);

lut_2_ro ro679(
   .en(en),
   .out(out[678]),
);

lut_2_ro ro680(
   .en(en),
   .out(out[679]),
);

lut_2_ro ro681(
   .en(en),
   .out(out[680]),
);

lut_2_ro ro682(
   .en(en),
   .out(out[681]),
);

lut_2_ro ro683(
   .en(en),
   .out(out[682]),
);

lut_2_ro ro684(
   .en(en),
   .out(out[683]),
);

lut_2_ro ro685(
   .en(en),
   .out(out[684]),
);

lut_2_ro ro686(
   .en(en),
   .out(out[685]),
);

lut_2_ro ro687(
   .en(en),
   .out(out[686]),
);

lut_2_ro ro688(
   .en(en),
   .out(out[687]),
);

lut_2_ro ro689(
   .en(en),
   .out(out[688]),
);

lut_2_ro ro690(
   .en(en),
   .out(out[689]),
);

lut_2_ro ro691(
   .en(en),
   .out(out[690]),
);

lut_2_ro ro692(
   .en(en),
   .out(out[691]),
);

lut_2_ro ro693(
   .en(en),
   .out(out[692]),
);

lut_2_ro ro694(
   .en(en),
   .out(out[693]),
);

lut_2_ro ro695(
   .en(en),
   .out(out[694]),
);

lut_2_ro ro696(
   .en(en),
   .out(out[695]),
);

lut_2_ro ro697(
   .en(en),
   .out(out[696]),
);

lut_2_ro ro698(
   .en(en),
   .out(out[697]),
);

lut_2_ro ro699(
   .en(en),
   .out(out[698]),
);

lut_2_ro ro700(
   .en(en),
   .out(out[699]),
);

lut_2_ro ro701(
   .en(en),
   .out(out[700]),
);

lut_2_ro ro702(
   .en(en),
   .out(out[701]),
);

lut_2_ro ro703(
   .en(en),
   .out(out[702]),
);

lut_2_ro ro704(
   .en(en),
   .out(out[703]),
);

lut_2_ro ro705(
   .en(en),
   .out(out[704]),
);

lut_2_ro ro706(
   .en(en),
   .out(out[705]),
);

lut_2_ro ro707(
   .en(en),
   .out(out[706]),
);

lut_2_ro ro708(
   .en(en),
   .out(out[707]),
);

lut_2_ro ro709(
   .en(en),
   .out(out[708]),
);

lut_2_ro ro710(
   .en(en),
   .out(out[709]),
);

lut_2_ro ro711(
   .en(en),
   .out(out[710]),
);

lut_2_ro ro712(
   .en(en),
   .out(out[711]),
);

lut_2_ro ro713(
   .en(en),
   .out(out[712]),
);

lut_2_ro ro714(
   .en(en),
   .out(out[713]),
);

lut_2_ro ro715(
   .en(en),
   .out(out[714]),
);

lut_2_ro ro716(
   .en(en),
   .out(out[715]),
);

lut_2_ro ro717(
   .en(en),
   .out(out[716]),
);

lut_2_ro ro718(
   .en(en),
   .out(out[717]),
);

lut_2_ro ro719(
   .en(en),
   .out(out[718]),
);

lut_2_ro ro720(
   .en(en),
   .out(out[719]),
);

lut_2_ro ro721(
   .en(en),
   .out(out[720]),
);

lut_2_ro ro722(
   .en(en),
   .out(out[721]),
);

lut_2_ro ro723(
   .en(en),
   .out(out[722]),
);

lut_2_ro ro724(
   .en(en),
   .out(out[723]),
);

lut_2_ro ro725(
   .en(en),
   .out(out[724]),
);

lut_2_ro ro726(
   .en(en),
   .out(out[725]),
);

lut_2_ro ro727(
   .en(en),
   .out(out[726]),
);

lut_2_ro ro728(
   .en(en),
   .out(out[727]),
);

lut_2_ro ro729(
   .en(en),
   .out(out[728]),
);

lut_2_ro ro730(
   .en(en),
   .out(out[729]),
);

lut_2_ro ro731(
   .en(en),
   .out(out[730]),
);

lut_2_ro ro732(
   .en(en),
   .out(out[731]),
);

lut_2_ro ro733(
   .en(en),
   .out(out[732]),
);

lut_2_ro ro734(
   .en(en),
   .out(out[733]),
);

lut_2_ro ro735(
   .en(en),
   .out(out[734]),
);

lut_2_ro ro736(
   .en(en),
   .out(out[735]),
);

lut_2_ro ro737(
   .en(en),
   .out(out[736]),
);

lut_2_ro ro738(
   .en(en),
   .out(out[737]),
);

lut_2_ro ro739(
   .en(en),
   .out(out[738]),
);

lut_2_ro ro740(
   .en(en),
   .out(out[739]),
);

lut_2_ro ro741(
   .en(en),
   .out(out[740]),
);

lut_2_ro ro742(
   .en(en),
   .out(out[741]),
);

lut_2_ro ro743(
   .en(en),
   .out(out[742]),
);

lut_2_ro ro744(
   .en(en),
   .out(out[743]),
);

lut_2_ro ro745(
   .en(en),
   .out(out[744]),
);

lut_2_ro ro746(
   .en(en),
   .out(out[745]),
);

lut_2_ro ro747(
   .en(en),
   .out(out[746]),
);

lut_2_ro ro748(
   .en(en),
   .out(out[747]),
);

lut_2_ro ro749(
   .en(en),
   .out(out[748]),
);

lut_2_ro ro750(
   .en(en),
   .out(out[749]),
);

lut_2_ro ro751(
   .en(en),
   .out(out[750]),
);

lut_2_ro ro752(
   .en(en),
   .out(out[751]),
);

lut_2_ro ro753(
   .en(en),
   .out(out[752]),
);

lut_2_ro ro754(
   .en(en),
   .out(out[753]),
);

lut_2_ro ro755(
   .en(en),
   .out(out[754]),
);

lut_2_ro ro756(
   .en(en),
   .out(out[755]),
);

lut_2_ro ro757(
   .en(en),
   .out(out[756]),
);

lut_2_ro ro758(
   .en(en),
   .out(out[757]),
);

lut_2_ro ro759(
   .en(en),
   .out(out[758]),
);

lut_2_ro ro760(
   .en(en),
   .out(out[759]),
);

lut_2_ro ro761(
   .en(en),
   .out(out[760]),
);

lut_2_ro ro762(
   .en(en),
   .out(out[761]),
);

lut_2_ro ro763(
   .en(en),
   .out(out[762]),
);

lut_2_ro ro764(
   .en(en),
   .out(out[763]),
);

lut_2_ro ro765(
   .en(en),
   .out(out[764]),
);

lut_2_ro ro766(
   .en(en),
   .out(out[765]),
);

lut_2_ro ro767(
   .en(en),
   .out(out[766]),
);

lut_2_ro ro768(
   .en(en),
   .out(out[767]),
);

lut_2_ro ro769(
   .en(en),
   .out(out[768]),
);

lut_2_ro ro770(
   .en(en),
   .out(out[769]),
);

lut_2_ro ro771(
   .en(en),
   .out(out[770]),
);

lut_2_ro ro772(
   .en(en),
   .out(out[771]),
);

lut_2_ro ro773(
   .en(en),
   .out(out[772]),
);

lut_2_ro ro774(
   .en(en),
   .out(out[773]),
);

lut_2_ro ro775(
   .en(en),
   .out(out[774]),
);

lut_2_ro ro776(
   .en(en),
   .out(out[775]),
);

lut_2_ro ro777(
   .en(en),
   .out(out[776]),
);

lut_2_ro ro778(
   .en(en),
   .out(out[777]),
);

lut_2_ro ro779(
   .en(en),
   .out(out[778]),
);

lut_2_ro ro780(
   .en(en),
   .out(out[779]),
);

lut_2_ro ro781(
   .en(en),
   .out(out[780]),
);

lut_2_ro ro782(
   .en(en),
   .out(out[781]),
);

lut_2_ro ro783(
   .en(en),
   .out(out[782]),
);

lut_2_ro ro784(
   .en(en),
   .out(out[783]),
);

lut_2_ro ro785(
   .en(en),
   .out(out[784]),
);

lut_2_ro ro786(
   .en(en),
   .out(out[785]),
);

lut_2_ro ro787(
   .en(en),
   .out(out[786]),
);

lut_2_ro ro788(
   .en(en),
   .out(out[787]),
);

lut_2_ro ro789(
   .en(en),
   .out(out[788]),
);

lut_2_ro ro790(
   .en(en),
   .out(out[789]),
);

lut_2_ro ro791(
   .en(en),
   .out(out[790]),
);

lut_2_ro ro792(
   .en(en),
   .out(out[791]),
);

lut_2_ro ro793(
   .en(en),
   .out(out[792]),
);

lut_2_ro ro794(
   .en(en),
   .out(out[793]),
);

lut_2_ro ro795(
   .en(en),
   .out(out[794]),
);

lut_2_ro ro796(
   .en(en),
   .out(out[795]),
);

lut_2_ro ro797(
   .en(en),
   .out(out[796]),
);

lut_2_ro ro798(
   .en(en),
   .out(out[797]),
);

lut_2_ro ro799(
   .en(en),
   .out(out[798]),
);

lut_2_ro ro800(
   .en(en),
   .out(out[799]),
);

lut_2_ro ro801(
   .en(en),
   .out(out[800]),
);

lut_2_ro ro802(
   .en(en),
   .out(out[801]),
);

lut_2_ro ro803(
   .en(en),
   .out(out[802]),
);

lut_2_ro ro804(
   .en(en),
   .out(out[803]),
);

lut_2_ro ro805(
   .en(en),
   .out(out[804]),
);

lut_2_ro ro806(
   .en(en),
   .out(out[805]),
);

lut_2_ro ro807(
   .en(en),
   .out(out[806]),
);

lut_2_ro ro808(
   .en(en),
   .out(out[807]),
);

lut_2_ro ro809(
   .en(en),
   .out(out[808]),
);

lut_2_ro ro810(
   .en(en),
   .out(out[809]),
);

lut_2_ro ro811(
   .en(en),
   .out(out[810]),
);

lut_2_ro ro812(
   .en(en),
   .out(out[811]),
);

lut_2_ro ro813(
   .en(en),
   .out(out[812]),
);

lut_2_ro ro814(
   .en(en),
   .out(out[813]),
);

lut_2_ro ro815(
   .en(en),
   .out(out[814]),
);

lut_2_ro ro816(
   .en(en),
   .out(out[815]),
);

lut_2_ro ro817(
   .en(en),
   .out(out[816]),
);

lut_2_ro ro818(
   .en(en),
   .out(out[817]),
);

lut_2_ro ro819(
   .en(en),
   .out(out[818]),
);

lut_2_ro ro820(
   .en(en),
   .out(out[819]),
);

lut_2_ro ro821(
   .en(en),
   .out(out[820]),
);

lut_2_ro ro822(
   .en(en),
   .out(out[821]),
);

lut_2_ro ro823(
   .en(en),
   .out(out[822]),
);

lut_2_ro ro824(
   .en(en),
   .out(out[823]),
);

lut_2_ro ro825(
   .en(en),
   .out(out[824]),
);

lut_2_ro ro826(
   .en(en),
   .out(out[825]),
);

lut_2_ro ro827(
   .en(en),
   .out(out[826]),
);

lut_2_ro ro828(
   .en(en),
   .out(out[827]),
);

lut_2_ro ro829(
   .en(en),
   .out(out[828]),
);

lut_2_ro ro830(
   .en(en),
   .out(out[829]),
);

lut_2_ro ro831(
   .en(en),
   .out(out[830]),
);

lut_2_ro ro832(
   .en(en),
   .out(out[831]),
);

lut_2_ro ro833(
   .en(en),
   .out(out[832]),
);

lut_2_ro ro834(
   .en(en),
   .out(out[833]),
);

lut_2_ro ro835(
   .en(en),
   .out(out[834]),
);

lut_2_ro ro836(
   .en(en),
   .out(out[835]),
);

lut_2_ro ro837(
   .en(en),
   .out(out[836]),
);

lut_2_ro ro838(
   .en(en),
   .out(out[837]),
);

lut_2_ro ro839(
   .en(en),
   .out(out[838]),
);

lut_2_ro ro840(
   .en(en),
   .out(out[839]),
);

lut_2_ro ro841(
   .en(en),
   .out(out[840]),
);

lut_2_ro ro842(
   .en(en),
   .out(out[841]),
);

lut_2_ro ro843(
   .en(en),
   .out(out[842]),
);

lut_2_ro ro844(
   .en(en),
   .out(out[843]),
);

lut_2_ro ro845(
   .en(en),
   .out(out[844]),
);

lut_2_ro ro846(
   .en(en),
   .out(out[845]),
);

lut_2_ro ro847(
   .en(en),
   .out(out[846]),
);

lut_2_ro ro848(
   .en(en),
   .out(out[847]),
);

lut_2_ro ro849(
   .en(en),
   .out(out[848]),
);

lut_2_ro ro850(
   .en(en),
   .out(out[849]),
);

lut_2_ro ro851(
   .en(en),
   .out(out[850]),
);

lut_2_ro ro852(
   .en(en),
   .out(out[851]),
);

lut_2_ro ro853(
   .en(en),
   .out(out[852]),
);

lut_2_ro ro854(
   .en(en),
   .out(out[853]),
);

lut_2_ro ro855(
   .en(en),
   .out(out[854]),
);

lut_2_ro ro856(
   .en(en),
   .out(out[855]),
);

lut_2_ro ro857(
   .en(en),
   .out(out[856]),
);

lut_2_ro ro858(
   .en(en),
   .out(out[857]),
);

lut_2_ro ro859(
   .en(en),
   .out(out[858]),
);

lut_2_ro ro860(
   .en(en),
   .out(out[859]),
);

lut_2_ro ro861(
   .en(en),
   .out(out[860]),
);

lut_2_ro ro862(
   .en(en),
   .out(out[861]),
);

lut_2_ro ro863(
   .en(en),
   .out(out[862]),
);

lut_2_ro ro864(
   .en(en),
   .out(out[863]),
);

lut_2_ro ro865(
   .en(en),
   .out(out[864]),
);

lut_2_ro ro866(
   .en(en),
   .out(out[865]),
);

lut_2_ro ro867(
   .en(en),
   .out(out[866]),
);

lut_2_ro ro868(
   .en(en),
   .out(out[867]),
);

lut_2_ro ro869(
   .en(en),
   .out(out[868]),
);

lut_2_ro ro870(
   .en(en),
   .out(out[869]),
);

lut_2_ro ro871(
   .en(en),
   .out(out[870]),
);

lut_2_ro ro872(
   .en(en),
   .out(out[871]),
);

lut_2_ro ro873(
   .en(en),
   .out(out[872]),
);

lut_2_ro ro874(
   .en(en),
   .out(out[873]),
);

lut_2_ro ro875(
   .en(en),
   .out(out[874]),
);

lut_2_ro ro876(
   .en(en),
   .out(out[875]),
);

lut_2_ro ro877(
   .en(en),
   .out(out[876]),
);

lut_2_ro ro878(
   .en(en),
   .out(out[877]),
);

lut_2_ro ro879(
   .en(en),
   .out(out[878]),
);

lut_2_ro ro880(
   .en(en),
   .out(out[879]),
);

lut_2_ro ro881(
   .en(en),
   .out(out[880]),
);

lut_2_ro ro882(
   .en(en),
   .out(out[881]),
);

lut_2_ro ro883(
   .en(en),
   .out(out[882]),
);

lut_2_ro ro884(
   .en(en),
   .out(out[883]),
);

lut_2_ro ro885(
   .en(en),
   .out(out[884]),
);

lut_2_ro ro886(
   .en(en),
   .out(out[885]),
);

lut_2_ro ro887(
   .en(en),
   .out(out[886]),
);

lut_2_ro ro888(
   .en(en),
   .out(out[887]),
);

lut_2_ro ro889(
   .en(en),
   .out(out[888]),
);

lut_2_ro ro890(
   .en(en),
   .out(out[889]),
);

lut_2_ro ro891(
   .en(en),
   .out(out[890]),
);

lut_2_ro ro892(
   .en(en),
   .out(out[891]),
);

lut_2_ro ro893(
   .en(en),
   .out(out[892]),
);

lut_2_ro ro894(
   .en(en),
   .out(out[893]),
);

lut_2_ro ro895(
   .en(en),
   .out(out[894]),
);

lut_2_ro ro896(
   .en(en),
   .out(out[895]),
);

lut_2_ro ro897(
   .en(en),
   .out(out[896]),
);

lut_2_ro ro898(
   .en(en),
   .out(out[897]),
);

lut_2_ro ro899(
   .en(en),
   .out(out[898]),
);

lut_2_ro ro900(
   .en(en),
   .out(out[899]),
);

lut_2_ro ro901(
   .en(en),
   .out(out[900]),
);

lut_2_ro ro902(
   .en(en),
   .out(out[901]),
);

lut_2_ro ro903(
   .en(en),
   .out(out[902]),
);

lut_2_ro ro904(
   .en(en),
   .out(out[903]),
);

lut_2_ro ro905(
   .en(en),
   .out(out[904]),
);

lut_2_ro ro906(
   .en(en),
   .out(out[905]),
);

lut_2_ro ro907(
   .en(en),
   .out(out[906]),
);

lut_2_ro ro908(
   .en(en),
   .out(out[907]),
);

lut_2_ro ro909(
   .en(en),
   .out(out[908]),
);

lut_2_ro ro910(
   .en(en),
   .out(out[909]),
);

lut_2_ro ro911(
   .en(en),
   .out(out[910]),
);

lut_2_ro ro912(
   .en(en),
   .out(out[911]),
);

lut_2_ro ro913(
   .en(en),
   .out(out[912]),
);

lut_2_ro ro914(
   .en(en),
   .out(out[913]),
);

lut_2_ro ro915(
   .en(en),
   .out(out[914]),
);

lut_2_ro ro916(
   .en(en),
   .out(out[915]),
);

lut_2_ro ro917(
   .en(en),
   .out(out[916]),
);

lut_2_ro ro918(
   .en(en),
   .out(out[917]),
);

lut_2_ro ro919(
   .en(en),
   .out(out[918]),
);

lut_2_ro ro920(
   .en(en),
   .out(out[919]),
);

lut_2_ro ro921(
   .en(en),
   .out(out[920]),
);

lut_2_ro ro922(
   .en(en),
   .out(out[921]),
);

lut_2_ro ro923(
   .en(en),
   .out(out[922]),
);

lut_2_ro ro924(
   .en(en),
   .out(out[923]),
);

lut_2_ro ro925(
   .en(en),
   .out(out[924]),
);

lut_2_ro ro926(
   .en(en),
   .out(out[925]),
);

lut_2_ro ro927(
   .en(en),
   .out(out[926]),
);

lut_2_ro ro928(
   .en(en),
   .out(out[927]),
);

lut_2_ro ro929(
   .en(en),
   .out(out[928]),
);

lut_2_ro ro930(
   .en(en),
   .out(out[929]),
);

lut_2_ro ro931(
   .en(en),
   .out(out[930]),
);

lut_2_ro ro932(
   .en(en),
   .out(out[931]),
);

lut_2_ro ro933(
   .en(en),
   .out(out[932]),
);

lut_2_ro ro934(
   .en(en),
   .out(out[933]),
);

lut_2_ro ro935(
   .en(en),
   .out(out[934]),
);

lut_2_ro ro936(
   .en(en),
   .out(out[935]),
);

lut_2_ro ro937(
   .en(en),
   .out(out[936]),
);

lut_2_ro ro938(
   .en(en),
   .out(out[937]),
);

lut_2_ro ro939(
   .en(en),
   .out(out[938]),
);

lut_2_ro ro940(
   .en(en),
   .out(out[939]),
);

lut_2_ro ro941(
   .en(en),
   .out(out[940]),
);

lut_2_ro ro942(
   .en(en),
   .out(out[941]),
);

lut_2_ro ro943(
   .en(en),
   .out(out[942]),
);

lut_2_ro ro944(
   .en(en),
   .out(out[943]),
);

lut_2_ro ro945(
   .en(en),
   .out(out[944]),
);

lut_2_ro ro946(
   .en(en),
   .out(out[945]),
);

lut_2_ro ro947(
   .en(en),
   .out(out[946]),
);

lut_2_ro ro948(
   .en(en),
   .out(out[947]),
);

lut_2_ro ro949(
   .en(en),
   .out(out[948]),
);

lut_2_ro ro950(
   .en(en),
   .out(out[949]),
);

lut_2_ro ro951(
   .en(en),
   .out(out[950]),
);

lut_2_ro ro952(
   .en(en),
   .out(out[951]),
);

lut_2_ro ro953(
   .en(en),
   .out(out[952]),
);

lut_2_ro ro954(
   .en(en),
   .out(out[953]),
);

lut_2_ro ro955(
   .en(en),
   .out(out[954]),
);

lut_2_ro ro956(
   .en(en),
   .out(out[955]),
);

lut_2_ro ro957(
   .en(en),
   .out(out[956]),
);

lut_2_ro ro958(
   .en(en),
   .out(out[957]),
);

lut_2_ro ro959(
   .en(en),
   .out(out[958]),
);

lut_2_ro ro960(
   .en(en),
   .out(out[959]),
);

lut_2_ro ro961(
   .en(en),
   .out(out[960]),
);

lut_2_ro ro962(
   .en(en),
   .out(out[961]),
);

lut_2_ro ro963(
   .en(en),
   .out(out[962]),
);

lut_2_ro ro964(
   .en(en),
   .out(out[963]),
);

lut_2_ro ro965(
   .en(en),
   .out(out[964]),
);

lut_2_ro ro966(
   .en(en),
   .out(out[965]),
);

lut_2_ro ro967(
   .en(en),
   .out(out[966]),
);

lut_2_ro ro968(
   .en(en),
   .out(out[967]),
);

lut_2_ro ro969(
   .en(en),
   .out(out[968]),
);

lut_2_ro ro970(
   .en(en),
   .out(out[969]),
);

lut_2_ro ro971(
   .en(en),
   .out(out[970]),
);

lut_2_ro ro972(
   .en(en),
   .out(out[971]),
);

lut_2_ro ro973(
   .en(en),
   .out(out[972]),
);

lut_2_ro ro974(
   .en(en),
   .out(out[973]),
);

lut_2_ro ro975(
   .en(en),
   .out(out[974]),
);

lut_2_ro ro976(
   .en(en),
   .out(out[975]),
);

lut_2_ro ro977(
   .en(en),
   .out(out[976]),
);

lut_2_ro ro978(
   .en(en),
   .out(out[977]),
);

lut_2_ro ro979(
   .en(en),
   .out(out[978]),
);

lut_2_ro ro980(
   .en(en),
   .out(out[979]),
);

lut_2_ro ro981(
   .en(en),
   .out(out[980]),
);

lut_2_ro ro982(
   .en(en),
   .out(out[981]),
);

lut_2_ro ro983(
   .en(en),
   .out(out[982]),
);

lut_2_ro ro984(
   .en(en),
   .out(out[983]),
);

lut_2_ro ro985(
   .en(en),
   .out(out[984]),
);

lut_2_ro ro986(
   .en(en),
   .out(out[985]),
);

lut_2_ro ro987(
   .en(en),
   .out(out[986]),
);

lut_2_ro ro988(
   .en(en),
   .out(out[987]),
);

lut_2_ro ro989(
   .en(en),
   .out(out[988]),
);

lut_2_ro ro990(
   .en(en),
   .out(out[989]),
);

lut_2_ro ro991(
   .en(en),
   .out(out[990]),
);

lut_2_ro ro992(
   .en(en),
   .out(out[991]),
);

lut_2_ro ro993(
   .en(en),
   .out(out[992]),
);

lut_2_ro ro994(
   .en(en),
   .out(out[993]),
);

lut_2_ro ro995(
   .en(en),
   .out(out[994]),
);

lut_2_ro ro996(
   .en(en),
   .out(out[995]),
);

lut_2_ro ro997(
   .en(en),
   .out(out[996]),
);

lut_2_ro ro998(
   .en(en),
   .out(out[997]),
);

lut_2_ro ro999(
   .en(en),
   .out(out[998]),
);

lut_2_ro ro1000(
   .en(en),
   .out(out[999]),
);

lut_2_ro ro1001(
   .en(en),
   .out(out[1000]),
);

lut_2_ro ro1002(
   .en(en),
   .out(out[1001]),
);

lut_2_ro ro1003(
   .en(en),
   .out(out[1002]),
);

lut_2_ro ro1004(
   .en(en),
   .out(out[1003]),
);

lut_2_ro ro1005(
   .en(en),
   .out(out[1004]),
);

lut_2_ro ro1006(
   .en(en),
   .out(out[1005]),
);

lut_2_ro ro1007(
   .en(en),
   .out(out[1006]),
);

lut_2_ro ro1008(
   .en(en),
   .out(out[1007]),
);

lut_2_ro ro1009(
   .en(en),
   .out(out[1008]),
);

lut_2_ro ro1010(
   .en(en),
   .out(out[1009]),
);

lut_2_ro ro1011(
   .en(en),
   .out(out[1010]),
);

lut_2_ro ro1012(
   .en(en),
   .out(out[1011]),
);

lut_2_ro ro1013(
   .en(en),
   .out(out[1012]),
);

lut_2_ro ro1014(
   .en(en),
   .out(out[1013]),
);

lut_2_ro ro1015(
   .en(en),
   .out(out[1014]),
);

lut_2_ro ro1016(
   .en(en),
   .out(out[1015]),
);

lut_2_ro ro1017(
   .en(en),
   .out(out[1016]),
);

lut_2_ro ro1018(
   .en(en),
   .out(out[1017]),
);

lut_2_ro ro1019(
   .en(en),
   .out(out[1018]),
);

lut_2_ro ro1020(
   .en(en),
   .out(out[1019]),
);

lut_2_ro ro1021(
   .en(en),
   .out(out[1020]),
);

lut_2_ro ro1022(
   .en(en),
   .out(out[1021]),
);

lut_2_ro ro1023(
   .en(en),
   .out(out[1022]),
);

lut_2_ro ro1024(
   .en(en),
   .out(out[1023]),
);

lut_2_ro ro1025(
   .en(en),
   .out(out[1024]),
);

lut_2_ro ro1026(
   .en(en),
   .out(out[1025]),
);

lut_2_ro ro1027(
   .en(en),
   .out(out[1026]),
);

lut_2_ro ro1028(
   .en(en),
   .out(out[1027]),
);

lut_2_ro ro1029(
   .en(en),
   .out(out[1028]),
);

lut_2_ro ro1030(
   .en(en),
   .out(out[1029]),
);

lut_2_ro ro1031(
   .en(en),
   .out(out[1030]),
);

lut_2_ro ro1032(
   .en(en),
   .out(out[1031]),
);

lut_2_ro ro1033(
   .en(en),
   .out(out[1032]),
);

lut_2_ro ro1034(
   .en(en),
   .out(out[1033]),
);

lut_2_ro ro1035(
   .en(en),
   .out(out[1034]),
);

lut_2_ro ro1036(
   .en(en),
   .out(out[1035]),
);

lut_2_ro ro1037(
   .en(en),
   .out(out[1036]),
);

lut_2_ro ro1038(
   .en(en),
   .out(out[1037]),
);

lut_2_ro ro1039(
   .en(en),
   .out(out[1038]),
);

lut_2_ro ro1040(
   .en(en),
   .out(out[1039]),
);

lut_2_ro ro1041(
   .en(en),
   .out(out[1040]),
);

lut_2_ro ro1042(
   .en(en),
   .out(out[1041]),
);

lut_2_ro ro1043(
   .en(en),
   .out(out[1042]),
);

lut_2_ro ro1044(
   .en(en),
   .out(out[1043]),
);

lut_2_ro ro1045(
   .en(en),
   .out(out[1044]),
);

lut_2_ro ro1046(
   .en(en),
   .out(out[1045]),
);

lut_2_ro ro1047(
   .en(en),
   .out(out[1046]),
);

lut_2_ro ro1048(
   .en(en),
   .out(out[1047]),
);

lut_2_ro ro1049(
   .en(en),
   .out(out[1048]),
);

lut_2_ro ro1050(
   .en(en),
   .out(out[1049]),
);

lut_2_ro ro1051(
   .en(en),
   .out(out[1050]),
);

lut_2_ro ro1052(
   .en(en),
   .out(out[1051]),
);

lut_2_ro ro1053(
   .en(en),
   .out(out[1052]),
);

lut_2_ro ro1054(
   .en(en),
   .out(out[1053]),
);

lut_2_ro ro1055(
   .en(en),
   .out(out[1054]),
);

lut_2_ro ro1056(
   .en(en),
   .out(out[1055]),
);

lut_2_ro ro1057(
   .en(en),
   .out(out[1056]),
);

lut_2_ro ro1058(
   .en(en),
   .out(out[1057]),
);

lut_2_ro ro1059(
   .en(en),
   .out(out[1058]),
);

lut_2_ro ro1060(
   .en(en),
   .out(out[1059]),
);

lut_2_ro ro1061(
   .en(en),
   .out(out[1060]),
);

lut_2_ro ro1062(
   .en(en),
   .out(out[1061]),
);

lut_2_ro ro1063(
   .en(en),
   .out(out[1062]),
);

lut_2_ro ro1064(
   .en(en),
   .out(out[1063]),
);

lut_2_ro ro1065(
   .en(en),
   .out(out[1064]),
);

lut_2_ro ro1066(
   .en(en),
   .out(out[1065]),
);

lut_2_ro ro1067(
   .en(en),
   .out(out[1066]),
);

lut_2_ro ro1068(
   .en(en),
   .out(out[1067]),
);

lut_2_ro ro1069(
   .en(en),
   .out(out[1068]),
);

lut_2_ro ro1070(
   .en(en),
   .out(out[1069]),
);

lut_2_ro ro1071(
   .en(en),
   .out(out[1070]),
);

lut_2_ro ro1072(
   .en(en),
   .out(out[1071]),
);

lut_2_ro ro1073(
   .en(en),
   .out(out[1072]),
);

lut_2_ro ro1074(
   .en(en),
   .out(out[1073]),
);

lut_2_ro ro1075(
   .en(en),
   .out(out[1074]),
);

lut_2_ro ro1076(
   .en(en),
   .out(out[1075]),
);

lut_2_ro ro1077(
   .en(en),
   .out(out[1076]),
);

lut_2_ro ro1078(
   .en(en),
   .out(out[1077]),
);

lut_2_ro ro1079(
   .en(en),
   .out(out[1078]),
);

lut_2_ro ro1080(
   .en(en),
   .out(out[1079]),
);

lut_2_ro ro1081(
   .en(en),
   .out(out[1080]),
);

lut_2_ro ro1082(
   .en(en),
   .out(out[1081]),
);

lut_2_ro ro1083(
   .en(en),
   .out(out[1082]),
);

lut_2_ro ro1084(
   .en(en),
   .out(out[1083]),
);

lut_2_ro ro1085(
   .en(en),
   .out(out[1084]),
);

lut_2_ro ro1086(
   .en(en),
   .out(out[1085]),
);

lut_2_ro ro1087(
   .en(en),
   .out(out[1086]),
);

lut_2_ro ro1088(
   .en(en),
   .out(out[1087]),
);

lut_2_ro ro1089(
   .en(en),
   .out(out[1088]),
);

lut_2_ro ro1090(
   .en(en),
   .out(out[1089]),
);

lut_2_ro ro1091(
   .en(en),
   .out(out[1090]),
);

lut_2_ro ro1092(
   .en(en),
   .out(out[1091]),
);

lut_2_ro ro1093(
   .en(en),
   .out(out[1092]),
);

lut_2_ro ro1094(
   .en(en),
   .out(out[1093]),
);

lut_2_ro ro1095(
   .en(en),
   .out(out[1094]),
);

lut_2_ro ro1096(
   .en(en),
   .out(out[1095]),
);

lut_2_ro ro1097(
   .en(en),
   .out(out[1096]),
);

lut_2_ro ro1098(
   .en(en),
   .out(out[1097]),
);

lut_2_ro ro1099(
   .en(en),
   .out(out[1098]),
);

lut_2_ro ro1100(
   .en(en),
   .out(out[1099]),
);
assign io_pad[13] = |out;
endmodule
