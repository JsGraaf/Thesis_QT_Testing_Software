
module MODULE_top(
   io_pad
);

// GPIO
inout    wire     [31:0]      io_pad      ;

assign io_pad[22] = io_pad[2];


(* keep = "true" *) wire lut_1_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut1 (
   .I0(io_pad[2]),
   .I1(lut_1_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_2_connect)
);

(* keep = "true" *) wire lut_2_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut2 (
   .I0(io_pad[2]),
   .I1(lut_2_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_3_connect)
);

(* keep = "true" *) wire lut_3_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut3 (
   .I0(io_pad[2]),
   .I1(lut_3_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_4_connect)
);

(* keep = "true" *) wire lut_4_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut4 (
   .I0(io_pad[2]),
   .I1(lut_4_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_5_connect)
);

(* keep = "true" *) wire lut_5_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut5 (
   .I0(io_pad[2]),
   .I1(lut_5_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_6_connect)
);

(* keep = "true" *) wire lut_6_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut6 (
   .I0(io_pad[2]),
   .I1(lut_6_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_7_connect)
);

(* keep = "true" *) wire lut_7_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut7 (
   .I0(io_pad[2]),
   .I1(lut_7_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_8_connect)
);

(* keep = "true" *) wire lut_8_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut8 (
   .I0(io_pad[2]),
   .I1(lut_8_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_9_connect)
);

(* keep = "true" *) wire lut_9_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut9 (
   .I0(io_pad[2]),
   .I1(lut_9_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_10_connect)
);

(* keep = "true" *) wire lut_10_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut10 (
   .I0(io_pad[2]),
   .I1(lut_10_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_11_connect)
);

(* keep = "true" *) wire lut_11_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut11 (
   .I0(io_pad[2]),
   .I1(lut_11_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_12_connect)
);

(* keep = "true" *) wire lut_12_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut12 (
   .I0(io_pad[2]),
   .I1(lut_12_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_13_connect)
);

(* keep = "true" *) wire lut_13_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut13 (
   .I0(io_pad[2]),
   .I1(lut_13_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_14_connect)
);

(* keep = "true" *) wire lut_14_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut14 (
   .I0(io_pad[2]),
   .I1(lut_14_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_15_connect)
);

(* keep = "true" *) wire lut_15_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut15 (
   .I0(io_pad[2]),
   .I1(lut_15_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_16_connect)
);

(* keep = "true" *) wire lut_16_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut16 (
   .I0(io_pad[2]),
   .I1(lut_16_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_17_connect)
);

(* keep = "true" *) wire lut_17_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut17 (
   .I0(io_pad[2]),
   .I1(lut_17_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_18_connect)
);

(* keep = "true" *) wire lut_18_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut18 (
   .I0(io_pad[2]),
   .I1(lut_18_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_19_connect)
);

(* keep = "true" *) wire lut_19_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut19 (
   .I0(io_pad[2]),
   .I1(lut_19_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_20_connect)
);

(* keep = "true" *) wire lut_20_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut20 (
   .I0(io_pad[2]),
   .I1(lut_20_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_21_connect)
);

(* keep = "true" *) wire lut_21_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut21 (
   .I0(io_pad[2]),
   .I1(lut_21_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_22_connect)
);

(* keep = "true" *) wire lut_22_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut22 (
   .I0(io_pad[2]),
   .I1(lut_22_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_23_connect)
);

(* keep = "true" *) wire lut_23_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut23 (
   .I0(io_pad[2]),
   .I1(lut_23_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_24_connect)
);

(* keep = "true" *) wire lut_24_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut24 (
   .I0(io_pad[2]),
   .I1(lut_24_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_25_connect)
);

(* keep = "true" *) wire lut_25_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut25 (
   .I0(io_pad[2]),
   .I1(lut_25_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_26_connect)
);

(* keep = "true" *) wire lut_26_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut26 (
   .I0(io_pad[2]),
   .I1(lut_26_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_27_connect)
);

(* keep = "true" *) wire lut_27_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut27 (
   .I0(io_pad[2]),
   .I1(lut_27_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_28_connect)
);

(* keep = "true" *) wire lut_28_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut28 (
   .I0(io_pad[2]),
   .I1(lut_28_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_29_connect)
);

(* keep = "true" *) wire lut_29_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut29 (
   .I0(io_pad[2]),
   .I1(lut_29_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_30_connect)
);

(* keep = "true" *) wire lut_30_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut30 (
   .I0(io_pad[2]),
   .I1(lut_30_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_31_connect)
);

(* keep = "true" *) wire lut_31_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut31 (
   .I0(io_pad[2]),
   .I1(lut_31_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_32_connect)
);

(* keep = "true" *) wire lut_32_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut32 (
   .I0(io_pad[2]),
   .I1(lut_32_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_33_connect)
);

(* keep = "true" *) wire lut_33_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut33 (
   .I0(io_pad[2]),
   .I1(lut_33_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_34_connect)
);

(* keep = "true" *) wire lut_34_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut34 (
   .I0(io_pad[2]),
   .I1(lut_34_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_35_connect)
);

(* keep = "true" *) wire lut_35_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut35 (
   .I0(io_pad[2]),
   .I1(lut_35_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_36_connect)
);

(* keep = "true" *) wire lut_36_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut36 (
   .I0(io_pad[2]),
   .I1(lut_36_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_37_connect)
);

(* keep = "true" *) wire lut_37_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut37 (
   .I0(io_pad[2]),
   .I1(lut_37_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_38_connect)
);

(* keep = "true" *) wire lut_38_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut38 (
   .I0(io_pad[2]),
   .I1(lut_38_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_39_connect)
);

(* keep = "true" *) wire lut_39_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut39 (
   .I0(io_pad[2]),
   .I1(lut_39_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_40_connect)
);

(* keep = "true" *) wire lut_40_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut40 (
   .I0(io_pad[2]),
   .I1(lut_40_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_41_connect)
);

(* keep = "true" *) wire lut_41_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut41 (
   .I0(io_pad[2]),
   .I1(lut_41_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_42_connect)
);

(* keep = "true" *) wire lut_42_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut42 (
   .I0(io_pad[2]),
   .I1(lut_42_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_43_connect)
);

(* keep = "true" *) wire lut_43_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut43 (
   .I0(io_pad[2]),
   .I1(lut_43_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_44_connect)
);

(* keep = "true" *) wire lut_44_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut44 (
   .I0(io_pad[2]),
   .I1(lut_44_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_45_connect)
);

(* keep = "true" *) wire lut_45_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut45 (
   .I0(io_pad[2]),
   .I1(lut_45_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_46_connect)
);

(* keep = "true" *) wire lut_46_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut46 (
   .I0(io_pad[2]),
   .I1(lut_46_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_47_connect)
);

(* keep = "true" *) wire lut_47_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut47 (
   .I0(io_pad[2]),
   .I1(lut_47_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_48_connect)
);

(* keep = "true" *) wire lut_48_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut48 (
   .I0(io_pad[2]),
   .I1(lut_48_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_49_connect)
);

(* keep = "true" *) wire lut_49_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut49 (
   .I0(io_pad[2]),
   .I1(lut_49_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_50_connect)
);

(* keep = "true" *) wire lut_50_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut50 (
   .I0(io_pad[2]),
   .I1(lut_50_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_51_connect)
);

(* keep = "true" *) wire lut_51_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut51 (
   .I0(io_pad[2]),
   .I1(lut_51_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_52_connect)
);

(* keep = "true" *) wire lut_52_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut52 (
   .I0(io_pad[2]),
   .I1(lut_52_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_53_connect)
);

(* keep = "true" *) wire lut_53_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut53 (
   .I0(io_pad[2]),
   .I1(lut_53_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_54_connect)
);

(* keep = "true" *) wire lut_54_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut54 (
   .I0(io_pad[2]),
   .I1(lut_54_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_55_connect)
);

(* keep = "true" *) wire lut_55_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut55 (
   .I0(io_pad[2]),
   .I1(lut_55_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_56_connect)
);

(* keep = "true" *) wire lut_56_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut56 (
   .I0(io_pad[2]),
   .I1(lut_56_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_57_connect)
);

(* keep = "true" *) wire lut_57_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut57 (
   .I0(io_pad[2]),
   .I1(lut_57_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_58_connect)
);

(* keep = "true" *) wire lut_58_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut58 (
   .I0(io_pad[2]),
   .I1(lut_58_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_59_connect)
);

(* keep = "true" *) wire lut_59_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut59 (
   .I0(io_pad[2]),
   .I1(lut_59_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_60_connect)
);

(* keep = "true" *) wire lut_60_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut60 (
   .I0(io_pad[2]),
   .I1(lut_60_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_61_connect)
);

(* keep = "true" *) wire lut_61_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut61 (
   .I0(io_pad[2]),
   .I1(lut_61_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_62_connect)
);

(* keep = "true" *) wire lut_62_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut62 (
   .I0(io_pad[2]),
   .I1(lut_62_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_63_connect)
);

(* keep = "true" *) wire lut_63_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut63 (
   .I0(io_pad[2]),
   .I1(lut_63_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_64_connect)
);

(* keep = "true" *) wire lut_64_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut64 (
   .I0(io_pad[2]),
   .I1(lut_64_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_65_connect)
);

(* keep = "true" *) wire lut_65_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut65 (
   .I0(io_pad[2]),
   .I1(lut_65_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_66_connect)
);

(* keep = "true" *) wire lut_66_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut66 (
   .I0(io_pad[2]),
   .I1(lut_66_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_67_connect)
);

(* keep = "true" *) wire lut_67_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut67 (
   .I0(io_pad[2]),
   .I1(lut_67_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_68_connect)
);

(* keep = "true" *) wire lut_68_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut68 (
   .I0(io_pad[2]),
   .I1(lut_68_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_69_connect)
);

(* keep = "true" *) wire lut_69_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut69 (
   .I0(io_pad[2]),
   .I1(lut_69_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_70_connect)
);

(* keep = "true" *) wire lut_70_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut70 (
   .I0(io_pad[2]),
   .I1(lut_70_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_71_connect)
);

(* keep = "true" *) wire lut_71_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut71 (
   .I0(io_pad[2]),
   .I1(lut_71_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_72_connect)
);

(* keep = "true" *) wire lut_72_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut72 (
   .I0(io_pad[2]),
   .I1(lut_72_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_73_connect)
);

(* keep = "true" *) wire lut_73_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut73 (
   .I0(io_pad[2]),
   .I1(lut_73_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_74_connect)
);

(* keep = "true" *) wire lut_74_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut74 (
   .I0(io_pad[2]),
   .I1(lut_74_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_75_connect)
);

(* keep = "true" *) wire lut_75_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut75 (
   .I0(io_pad[2]),
   .I1(lut_75_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_76_connect)
);

(* keep = "true" *) wire lut_76_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut76 (
   .I0(io_pad[2]),
   .I1(lut_76_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_77_connect)
);

(* keep = "true" *) wire lut_77_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut77 (
   .I0(io_pad[2]),
   .I1(lut_77_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_78_connect)
);

(* keep = "true" *) wire lut_78_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut78 (
   .I0(io_pad[2]),
   .I1(lut_78_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_79_connect)
);

(* keep = "true" *) wire lut_79_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut79 (
   .I0(io_pad[2]),
   .I1(lut_79_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_80_connect)
);

(* keep = "true" *) wire lut_80_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut80 (
   .I0(io_pad[2]),
   .I1(lut_80_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_81_connect)
);

(* keep = "true" *) wire lut_81_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut81 (
   .I0(io_pad[2]),
   .I1(lut_81_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_82_connect)
);

(* keep = "true" *) wire lut_82_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut82 (
   .I0(io_pad[2]),
   .I1(lut_82_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_83_connect)
);

(* keep = "true" *) wire lut_83_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut83 (
   .I0(io_pad[2]),
   .I1(lut_83_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_84_connect)
);

(* keep = "true" *) wire lut_84_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut84 (
   .I0(io_pad[2]),
   .I1(lut_84_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_85_connect)
);

(* keep = "true" *) wire lut_85_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut85 (
   .I0(io_pad[2]),
   .I1(lut_85_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_86_connect)
);

(* keep = "true" *) wire lut_86_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut86 (
   .I0(io_pad[2]),
   .I1(lut_86_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_87_connect)
);

(* keep = "true" *) wire lut_87_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut87 (
   .I0(io_pad[2]),
   .I1(lut_87_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_88_connect)
);

(* keep = "true" *) wire lut_88_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut88 (
   .I0(io_pad[2]),
   .I1(lut_88_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_89_connect)
);

(* keep = "true" *) wire lut_89_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut89 (
   .I0(io_pad[2]),
   .I1(lut_89_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_90_connect)
);

(* keep = "true" *) wire lut_90_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut90 (
   .I0(io_pad[2]),
   .I1(lut_90_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_91_connect)
);

(* keep = "true" *) wire lut_91_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut91 (
   .I0(io_pad[2]),
   .I1(lut_91_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_92_connect)
);

(* keep = "true" *) wire lut_92_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut92 (
   .I0(io_pad[2]),
   .I1(lut_92_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_93_connect)
);

(* keep = "true" *) wire lut_93_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut93 (
   .I0(io_pad[2]),
   .I1(lut_93_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_94_connect)
);

(* keep = "true" *) wire lut_94_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut94 (
   .I0(io_pad[2]),
   .I1(lut_94_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_95_connect)
);

(* keep = "true" *) wire lut_95_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut95 (
   .I0(io_pad[2]),
   .I1(lut_95_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_96_connect)
);

(* keep = "true" *) wire lut_96_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut96 (
   .I0(io_pad[2]),
   .I1(lut_96_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_97_connect)
);

(* keep = "true" *) wire lut_97_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut97 (
   .I0(io_pad[2]),
   .I1(lut_97_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_98_connect)
);

(* keep = "true" *) wire lut_98_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut98 (
   .I0(io_pad[2]),
   .I1(lut_98_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_99_connect)
);

(* keep = "true" *) wire lut_99_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut99 (
   .I0(io_pad[2]),
   .I1(lut_99_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_100_connect)
);

(* keep = "true" *) wire lut_100_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut100 (
   .I0(io_pad[2]),
   .I1(lut_100_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_101_connect)
);

(* keep = "true" *) wire lut_101_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut101 (
   .I0(io_pad[2]),
   .I1(lut_101_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_102_connect)
);

(* keep = "true" *) wire lut_102_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut102 (
   .I0(io_pad[2]),
   .I1(lut_102_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_103_connect)
);

(* keep = "true" *) wire lut_103_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut103 (
   .I0(io_pad[2]),
   .I1(lut_103_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_104_connect)
);

(* keep = "true" *) wire lut_104_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut104 (
   .I0(io_pad[2]),
   .I1(lut_104_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_105_connect)
);

(* keep = "true" *) wire lut_105_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut105 (
   .I0(io_pad[2]),
   .I1(lut_105_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_106_connect)
);

(* keep = "true" *) wire lut_106_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut106 (
   .I0(io_pad[2]),
   .I1(lut_106_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_107_connect)
);

(* keep = "true" *) wire lut_107_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut107 (
   .I0(io_pad[2]),
   .I1(lut_107_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_108_connect)
);

(* keep = "true" *) wire lut_108_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut108 (
   .I0(io_pad[2]),
   .I1(lut_108_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_109_connect)
);

(* keep = "true" *) wire lut_109_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut109 (
   .I0(io_pad[2]),
   .I1(lut_109_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_110_connect)
);

(* keep = "true" *) wire lut_110_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut110 (
   .I0(io_pad[2]),
   .I1(lut_110_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_111_connect)
);

(* keep = "true" *) wire lut_111_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut111 (
   .I0(io_pad[2]),
   .I1(lut_111_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_112_connect)
);

(* keep = "true" *) wire lut_112_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut112 (
   .I0(io_pad[2]),
   .I1(lut_112_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_113_connect)
);

(* keep = "true" *) wire lut_113_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut113 (
   .I0(io_pad[2]),
   .I1(lut_113_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_114_connect)
);

(* keep = "true" *) wire lut_114_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut114 (
   .I0(io_pad[2]),
   .I1(lut_114_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_115_connect)
);

(* keep = "true" *) wire lut_115_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut115 (
   .I0(io_pad[2]),
   .I1(lut_115_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_116_connect)
);

(* keep = "true" *) wire lut_116_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut116 (
   .I0(io_pad[2]),
   .I1(lut_116_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_117_connect)
);

(* keep = "true" *) wire lut_117_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut117 (
   .I0(io_pad[2]),
   .I1(lut_117_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_118_connect)
);

(* keep = "true" *) wire lut_118_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut118 (
   .I0(io_pad[2]),
   .I1(lut_118_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_119_connect)
);

(* keep = "true" *) wire lut_119_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut119 (
   .I0(io_pad[2]),
   .I1(lut_119_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_120_connect)
);

(* keep = "true" *) wire lut_120_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut120 (
   .I0(io_pad[2]),
   .I1(lut_120_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_121_connect)
);

(* keep = "true" *) wire lut_121_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut121 (
   .I0(io_pad[2]),
   .I1(lut_121_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_122_connect)
);

(* keep = "true" *) wire lut_122_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut122 (
   .I0(io_pad[2]),
   .I1(lut_122_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_123_connect)
);

(* keep = "true" *) wire lut_123_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut123 (
   .I0(io_pad[2]),
   .I1(lut_123_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_124_connect)
);

(* keep = "true" *) wire lut_124_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut124 (
   .I0(io_pad[2]),
   .I1(lut_124_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_125_connect)
);

(* keep = "true" *) wire lut_125_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut125 (
   .I0(io_pad[2]),
   .I1(lut_125_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_126_connect)
);

(* keep = "true" *) wire lut_126_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut126 (
   .I0(io_pad[2]),
   .I1(lut_126_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_127_connect)
);

(* keep = "true" *) wire lut_127_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut127 (
   .I0(io_pad[2]),
   .I1(lut_127_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_128_connect)
);

(* keep = "true" *) wire lut_128_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut128 (
   .I0(io_pad[2]),
   .I1(lut_128_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_129_connect)
);

(* keep = "true" *) wire lut_129_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut129 (
   .I0(io_pad[2]),
   .I1(lut_129_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_130_connect)
);

(* keep = "true" *) wire lut_130_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut130 (
   .I0(io_pad[2]),
   .I1(lut_130_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_131_connect)
);

(* keep = "true" *) wire lut_131_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut131 (
   .I0(io_pad[2]),
   .I1(lut_131_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_132_connect)
);

(* keep = "true" *) wire lut_132_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut132 (
   .I0(io_pad[2]),
   .I1(lut_132_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_133_connect)
);

(* keep = "true" *) wire lut_133_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut133 (
   .I0(io_pad[2]),
   .I1(lut_133_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_134_connect)
);

(* keep = "true" *) wire lut_134_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut134 (
   .I0(io_pad[2]),
   .I1(lut_134_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_135_connect)
);

(* keep = "true" *) wire lut_135_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut135 (
   .I0(io_pad[2]),
   .I1(lut_135_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_136_connect)
);

(* keep = "true" *) wire lut_136_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut136 (
   .I0(io_pad[2]),
   .I1(lut_136_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_137_connect)
);

(* keep = "true" *) wire lut_137_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut137 (
   .I0(io_pad[2]),
   .I1(lut_137_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_138_connect)
);

(* keep = "true" *) wire lut_138_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut138 (
   .I0(io_pad[2]),
   .I1(lut_138_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_139_connect)
);

(* keep = "true" *) wire lut_139_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut139 (
   .I0(io_pad[2]),
   .I1(lut_139_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_140_connect)
);

(* keep = "true" *) wire lut_140_connect;
(* keep = "true" *) LUT4 #(
   .INIT(16'b0000000000000010)
) lut140 (
   .I0(io_pad[2]),
   .I1(lut_140_connect),
   .I2(1'b0),
   .I3(1'b0),
   .O(lut_141_connect)
);
endmodule
