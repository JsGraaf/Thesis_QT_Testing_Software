
module MODULE_top(
   io_pad
);

// GPIO
inout       wire    [31:0]      io_pad          ;

wire connectWire0;
assign io_pad[6] = connectWire0; 

wire connectWire1;
inv invert1 (
   .A(connectWire0),
   .Q(connectWire1)
);

wire connectWire2;
inv invert2 (
   .A(connectWire1),
   .Q(connectWire2)
);

wire connectWire3;
inv invert3 (
   .A(connectWire2),
   .Q(connectWire3)
);

wire connectWire4;
inv invert4 (
   .A(connectWire3),
   .Q(connectWire4)
);

wire connectWire5;
inv invert5 (
   .A(connectWire4),
   .Q(connectWire5)
);

wire connectWire6;
inv invert6 (
   .A(connectWire5),
   .Q(connectWire6)
);

wire connectWire7;
inv invert7 (
   .A(connectWire6),
   .Q(connectWire7)
);

wire connectWire8;
inv invert8 (
   .A(connectWire7),
   .Q(connectWire8)
);

wire connectWire9;
inv invert9 (
   .A(connectWire8),
   .Q(connectWire9)
);

wire connectWire10;
inv invert10 (
   .A(connectWire9),
   .Q(connectWire10)
);

wire connectWire11;
inv invert11 (
   .A(connectWire10),
   .Q(connectWire11)
);

wire connectWire12;
inv invert12 (
   .A(connectWire11),
   .Q(connectWire12)
);

wire connectWire13;
inv invert13 (
   .A(connectWire12),
   .Q(connectWire13)
);

wire connectWire14;
inv invert14 (
   .A(connectWire13),
   .Q(connectWire14)
);

wire connectWire15;
inv invert15 (
   .A(connectWire14),
   .Q(connectWire15)
);

wire connectWire16;
inv invert16 (
   .A(connectWire15),
   .Q(connectWire16)
);

wire connectWire17;
inv invert17 (
   .A(connectWire16),
   .Q(connectWire17)
);

wire connectWire18;
inv invert18 (
   .A(connectWire17),
   .Q(connectWire18)
);

wire connectWire19;
inv invert19 (
   .A(connectWire18),
   .Q(connectWire19)
);

wire connectWire20;
inv invert20 (
   .A(connectWire19),
   .Q(connectWire20)
);

wire connectWire21;
inv invert21 (
   .A(connectWire20),
   .Q(connectWire21)
);

wire connectWire22;
inv invert22 (
   .A(connectWire21),
   .Q(connectWire22)
);

wire connectWire23;
inv invert23 (
   .A(connectWire22),
   .Q(connectWire23)
);

wire connectWire24;
inv invert24 (
   .A(connectWire23),
   .Q(connectWire24)
);

wire connectWire25;
inv invert25 (
   .A(connectWire24),
   .Q(connectWire25)
);

wire connectWire26;
inv invert26 (
   .A(connectWire25),
   .Q(connectWire26)
);

wire connectWire27;
inv invert27 (
   .A(connectWire26),
   .Q(connectWire27)
);

wire connectWire28;
inv invert28 (
   .A(connectWire27),
   .Q(connectWire28)
);

wire connectWire29;
inv invert29 (
   .A(connectWire28),
   .Q(connectWire29)
);

wire connectWire30;
inv invert30 (
   .A(connectWire29),
   .Q(connectWire30)
);

wire connectWire31;
inv invert31 (
   .A(connectWire30),
   .Q(connectWire31)
);

wire connectWire32;
inv invert32 (
   .A(connectWire31),
   .Q(connectWire32)
);

wire connectWire33;
inv invert33 (
   .A(connectWire32),
   .Q(connectWire33)
);

wire connectWire34;
inv invert34 (
   .A(connectWire33),
   .Q(connectWire34)
);

wire connectWire35;
inv invert35 (
   .A(connectWire34),
   .Q(connectWire35)
);

wire connectWire36;
inv invert36 (
   .A(connectWire35),
   .Q(connectWire36)
);

wire connectWire37;
inv invert37 (
   .A(connectWire36),
   .Q(connectWire37)
);

wire connectWire38;
inv invert38 (
   .A(connectWire37),
   .Q(connectWire38)
);

wire connectWire39;
inv invert39 (
   .A(connectWire38),
   .Q(connectWire39)
);

wire connectWire40;
inv invert40 (
   .A(connectWire39),
   .Q(connectWire40)
);

wire connectWire41;
inv invert41 (
   .A(connectWire40),
   .Q(connectWire41)
);

wire connectWire42;
inv invert42 (
   .A(connectWire41),
   .Q(connectWire42)
);

wire connectWire43;
inv invert43 (
   .A(connectWire42),
   .Q(connectWire43)
);

wire connectWire44;
inv invert44 (
   .A(connectWire43),
   .Q(connectWire44)
);

wire connectWire45;
inv invert45 (
   .A(connectWire44),
   .Q(connectWire45)
);

wire connectWire46;
inv invert46 (
   .A(connectWire45),
   .Q(connectWire46)
);

wire connectWire47;
inv invert47 (
   .A(connectWire46),
   .Q(connectWire47)
);

wire connectWire48;
inv invert48 (
   .A(connectWire47),
   .Q(connectWire48)
);

wire connectWire49;
inv invert49 (
   .A(connectWire48),
   .Q(connectWire49)
);

wire connectWire50;
inv invert50 (
   .A(connectWire49),
   .Q(connectWire50)
);

wire connectWire51;
inv invert51 (
   .A(connectWire50),
   .Q(connectWire51)
);

wire connectWire52;
inv invert52 (
   .A(connectWire51),
   .Q(connectWire52)
);

wire connectWire53;
inv invert53 (
   .A(connectWire52),
   .Q(connectWire53)
);

wire connectWire54;
inv invert54 (
   .A(connectWire53),
   .Q(connectWire54)
);

wire connectWire55;
inv invert55 (
   .A(connectWire54),
   .Q(connectWire55)
);

wire connectWire56;
inv invert56 (
   .A(connectWire55),
   .Q(connectWire56)
);

wire connectWire57;
inv invert57 (
   .A(connectWire56),
   .Q(connectWire57)
);

wire connectWire58;
inv invert58 (
   .A(connectWire57),
   .Q(connectWire58)
);

wire connectWire59;
inv invert59 (
   .A(connectWire58),
   .Q(connectWire59)
);

wire connectWire60;
inv invert60 (
   .A(connectWire59),
   .Q(connectWire60)
);

wire connectWire61;
inv invert61 (
   .A(connectWire60),
   .Q(connectWire61)
);

wire connectWire62;
inv invert62 (
   .A(connectWire61),
   .Q(connectWire62)
);

wire connectWire63;
inv invert63 (
   .A(connectWire62),
   .Q(connectWire63)
);

wire connectWire64;
inv invert64 (
   .A(connectWire63),
   .Q(connectWire64)
);

wire connectWire65;
inv invert65 (
   .A(connectWire64),
   .Q(connectWire65)
);

wire connectWire66;
inv invert66 (
   .A(connectWire65),
   .Q(connectWire66)
);

wire connectWire67;
inv invert67 (
   .A(connectWire66),
   .Q(connectWire67)
);

wire connectWire68;
inv invert68 (
   .A(connectWire67),
   .Q(connectWire68)
);

wire connectWire69;
inv invert69 (
   .A(connectWire68),
   .Q(connectWire69)
);

wire connectWire70;
inv invert70 (
   .A(connectWire69),
   .Q(connectWire70)
);

assign io_pad[21] = connectWire70;
endmodule
