module mux8_ro(
   input en,
   output out,
);

(*keep*)wire connect;

assign connect = en ? connect : 0;
assign out = en ? connect : 0;

mux8x0 ro (
   .S0(connect),
   .S1(1'b0),
   .S2(1'b0),
   .A(1'b1),
   .B(1'b0),
   .C(1'b0),
   .D(1'b0),
   .E(1'b0),
   .F(1'b0),
   .G(1'b0),
   .H(1'b0),
   .Q(connect)
);
endmodule

 
module MODULE_top(
   io_pad
);

// GPIO
inout    wire     [31:0]      io_pad      ;

wire [149:0] out;

reg en;
initial begin
   en <= 1;
end

mux8_ro ro1(
   .en(en),
   .out(out[0]),
);

mux8_ro ro2(
   .en(en),
   .out(out[1]),
);

mux8_ro ro3(
   .en(en),
   .out(out[2]),
);

mux8_ro ro4(
   .en(en),
   .out(out[3]),
);

mux8_ro ro5(
   .en(en),
   .out(out[4]),
);

mux8_ro ro6(
   .en(en),
   .out(out[5]),
);

mux8_ro ro7(
   .en(en),
   .out(out[6]),
);

mux8_ro ro8(
   .en(en),
   .out(out[7]),
);

mux8_ro ro9(
   .en(en),
   .out(out[8]),
);

mux8_ro ro10(
   .en(en),
   .out(out[9]),
);

mux8_ro ro11(
   .en(en),
   .out(out[10]),
);

mux8_ro ro12(
   .en(en),
   .out(out[11]),
);

mux8_ro ro13(
   .en(en),
   .out(out[12]),
);

mux8_ro ro14(
   .en(en),
   .out(out[13]),
);

mux8_ro ro15(
   .en(en),
   .out(out[14]),
);

mux8_ro ro16(
   .en(en),
   .out(out[15]),
);

mux8_ro ro17(
   .en(en),
   .out(out[16]),
);

mux8_ro ro18(
   .en(en),
   .out(out[17]),
);

mux8_ro ro19(
   .en(en),
   .out(out[18]),
);

mux8_ro ro20(
   .en(en),
   .out(out[19]),
);

mux8_ro ro21(
   .en(en),
   .out(out[20]),
);

mux8_ro ro22(
   .en(en),
   .out(out[21]),
);

mux8_ro ro23(
   .en(en),
   .out(out[22]),
);

mux8_ro ro24(
   .en(en),
   .out(out[23]),
);

mux8_ro ro25(
   .en(en),
   .out(out[24]),
);

mux8_ro ro26(
   .en(en),
   .out(out[25]),
);

mux8_ro ro27(
   .en(en),
   .out(out[26]),
);

mux8_ro ro28(
   .en(en),
   .out(out[27]),
);

mux8_ro ro29(
   .en(en),
   .out(out[28]),
);

mux8_ro ro30(
   .en(en),
   .out(out[29]),
);

mux8_ro ro31(
   .en(en),
   .out(out[30]),
);

mux8_ro ro32(
   .en(en),
   .out(out[31]),
);

mux8_ro ro33(
   .en(en),
   .out(out[32]),
);

mux8_ro ro34(
   .en(en),
   .out(out[33]),
);

mux8_ro ro35(
   .en(en),
   .out(out[34]),
);

mux8_ro ro36(
   .en(en),
   .out(out[35]),
);

mux8_ro ro37(
   .en(en),
   .out(out[36]),
);

mux8_ro ro38(
   .en(en),
   .out(out[37]),
);

mux8_ro ro39(
   .en(en),
   .out(out[38]),
);

mux8_ro ro40(
   .en(en),
   .out(out[39]),
);

mux8_ro ro41(
   .en(en),
   .out(out[40]),
);

mux8_ro ro42(
   .en(en),
   .out(out[41]),
);

mux8_ro ro43(
   .en(en),
   .out(out[42]),
);

mux8_ro ro44(
   .en(en),
   .out(out[43]),
);

mux8_ro ro45(
   .en(en),
   .out(out[44]),
);

mux8_ro ro46(
   .en(en),
   .out(out[45]),
);

mux8_ro ro47(
   .en(en),
   .out(out[46]),
);

mux8_ro ro48(
   .en(en),
   .out(out[47]),
);

mux8_ro ro49(
   .en(en),
   .out(out[48]),
);

mux8_ro ro50(
   .en(en),
   .out(out[49]),
);

mux8_ro ro51(
   .en(en),
   .out(out[50]),
);

mux8_ro ro52(
   .en(en),
   .out(out[51]),
);

mux8_ro ro53(
   .en(en),
   .out(out[52]),
);

mux8_ro ro54(
   .en(en),
   .out(out[53]),
);

mux8_ro ro55(
   .en(en),
   .out(out[54]),
);

mux8_ro ro56(
   .en(en),
   .out(out[55]),
);

mux8_ro ro57(
   .en(en),
   .out(out[56]),
);

mux8_ro ro58(
   .en(en),
   .out(out[57]),
);

mux8_ro ro59(
   .en(en),
   .out(out[58]),
);

mux8_ro ro60(
   .en(en),
   .out(out[59]),
);

mux8_ro ro61(
   .en(en),
   .out(out[60]),
);

mux8_ro ro62(
   .en(en),
   .out(out[61]),
);

mux8_ro ro63(
   .en(en),
   .out(out[62]),
);

mux8_ro ro64(
   .en(en),
   .out(out[63]),
);

mux8_ro ro65(
   .en(en),
   .out(out[64]),
);

mux8_ro ro66(
   .en(en),
   .out(out[65]),
);

mux8_ro ro67(
   .en(en),
   .out(out[66]),
);

mux8_ro ro68(
   .en(en),
   .out(out[67]),
);

mux8_ro ro69(
   .en(en),
   .out(out[68]),
);

mux8_ro ro70(
   .en(en),
   .out(out[69]),
);

mux8_ro ro71(
   .en(en),
   .out(out[70]),
);

mux8_ro ro72(
   .en(en),
   .out(out[71]),
);

mux8_ro ro73(
   .en(en),
   .out(out[72]),
);

mux8_ro ro74(
   .en(en),
   .out(out[73]),
);

mux8_ro ro75(
   .en(en),
   .out(out[74]),
);

mux8_ro ro76(
   .en(en),
   .out(out[75]),
);

mux8_ro ro77(
   .en(en),
   .out(out[76]),
);

mux8_ro ro78(
   .en(en),
   .out(out[77]),
);

mux8_ro ro79(
   .en(en),
   .out(out[78]),
);

mux8_ro ro80(
   .en(en),
   .out(out[79]),
);

mux8_ro ro81(
   .en(en),
   .out(out[80]),
);

mux8_ro ro82(
   .en(en),
   .out(out[81]),
);

mux8_ro ro83(
   .en(en),
   .out(out[82]),
);

mux8_ro ro84(
   .en(en),
   .out(out[83]),
);

mux8_ro ro85(
   .en(en),
   .out(out[84]),
);

mux8_ro ro86(
   .en(en),
   .out(out[85]),
);

mux8_ro ro87(
   .en(en),
   .out(out[86]),
);

mux8_ro ro88(
   .en(en),
   .out(out[87]),
);

mux8_ro ro89(
   .en(en),
   .out(out[88]),
);

mux8_ro ro90(
   .en(en),
   .out(out[89]),
);

mux8_ro ro91(
   .en(en),
   .out(out[90]),
);

mux8_ro ro92(
   .en(en),
   .out(out[91]),
);

mux8_ro ro93(
   .en(en),
   .out(out[92]),
);

mux8_ro ro94(
   .en(en),
   .out(out[93]),
);

mux8_ro ro95(
   .en(en),
   .out(out[94]),
);

mux8_ro ro96(
   .en(en),
   .out(out[95]),
);

mux8_ro ro97(
   .en(en),
   .out(out[96]),
);

mux8_ro ro98(
   .en(en),
   .out(out[97]),
);

mux8_ro ro99(
   .en(en),
   .out(out[98]),
);

mux8_ro ro100(
   .en(en),
   .out(out[99]),
);

mux8_ro ro101(
   .en(en),
   .out(out[100]),
);

mux8_ro ro102(
   .en(en),
   .out(out[101]),
);

mux8_ro ro103(
   .en(en),
   .out(out[102]),
);

mux8_ro ro104(
   .en(en),
   .out(out[103]),
);

mux8_ro ro105(
   .en(en),
   .out(out[104]),
);

mux8_ro ro106(
   .en(en),
   .out(out[105]),
);

mux8_ro ro107(
   .en(en),
   .out(out[106]),
);

mux8_ro ro108(
   .en(en),
   .out(out[107]),
);

mux8_ro ro109(
   .en(en),
   .out(out[108]),
);

mux8_ro ro110(
   .en(en),
   .out(out[109]),
);

mux8_ro ro111(
   .en(en),
   .out(out[110]),
);

mux8_ro ro112(
   .en(en),
   .out(out[111]),
);

mux8_ro ro113(
   .en(en),
   .out(out[112]),
);

mux8_ro ro114(
   .en(en),
   .out(out[113]),
);

mux8_ro ro115(
   .en(en),
   .out(out[114]),
);

mux8_ro ro116(
   .en(en),
   .out(out[115]),
);

mux8_ro ro117(
   .en(en),
   .out(out[116]),
);

mux8_ro ro118(
   .en(en),
   .out(out[117]),
);

mux8_ro ro119(
   .en(en),
   .out(out[118]),
);

mux8_ro ro120(
   .en(en),
   .out(out[119]),
);

mux8_ro ro121(
   .en(en),
   .out(out[120]),
);

mux8_ro ro122(
   .en(en),
   .out(out[121]),
);

mux8_ro ro123(
   .en(en),
   .out(out[122]),
);

mux8_ro ro124(
   .en(en),
   .out(out[123]),
);

mux8_ro ro125(
   .en(en),
   .out(out[124]),
);

mux8_ro ro126(
   .en(en),
   .out(out[125]),
);

mux8_ro ro127(
   .en(en),
   .out(out[126]),
);

mux8_ro ro128(
   .en(en),
   .out(out[127]),
);

mux8_ro ro129(
   .en(en),
   .out(out[128]),
);

mux8_ro ro130(
   .en(en),
   .out(out[129]),
);

mux8_ro ro131(
   .en(en),
   .out(out[130]),
);

mux8_ro ro132(
   .en(en),
   .out(out[131]),
);

mux8_ro ro133(
   .en(en),
   .out(out[132]),
);

mux8_ro ro134(
   .en(en),
   .out(out[133]),
);

mux8_ro ro135(
   .en(en),
   .out(out[134]),
);

mux8_ro ro136(
   .en(en),
   .out(out[135]),
);

mux8_ro ro137(
   .en(en),
   .out(out[136]),
);

mux8_ro ro138(
   .en(en),
   .out(out[137]),
);

mux8_ro ro139(
   .en(en),
   .out(out[138]),
);

mux8_ro ro140(
   .en(en),
   .out(out[139]),
);

mux8_ro ro141(
   .en(en),
   .out(out[140]),
);

mux8_ro ro142(
   .en(en),
   .out(out[141]),
);

mux8_ro ro143(
   .en(en),
   .out(out[142]),
);

mux8_ro ro144(
   .en(en),
   .out(out[143]),
);

mux8_ro ro145(
   .en(en),
   .out(out[144]),
);

mux8_ro ro146(
   .en(en),
   .out(out[145]),
);

mux8_ro ro147(
   .en(en),
   .out(out[146]),
);

mux8_ro ro148(
   .en(en),
   .out(out[147]),
);

mux8_ro ro149(
   .en(en),
   .out(out[148]),
);

mux8_ro ro150(
   .en(en),
   .out(out[149]),
);

assign io_pad[13] = |out;
endmodule
