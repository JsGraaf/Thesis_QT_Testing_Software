module not_3_ro(
   input en,
   output out,
);

assign connect[0] = en ? connect[3] : 0;
assign out = en ? connect[3] : 0;

(*keep*)wire [3:0] connect;

inv inv1 (
   .A(connect[0]),
   .Q(connect[1])
);

inv inv2 (
   .A(connect[1]),
   .Q(connect[2]),
);

inv inv3 (
   .A(connect[2]),
   .Q(connect[3])
);
endmodule

module MODULE_top(
   io_pad
);

// GPIO
inout    wire     [31:0]      io_pad      ;

wire [189:0] out;

reg en;
initial begin
   en <= 1;
end

not_3_ro ro0 (
   .en(en),
   .out(out[0]),
);

not_3_ro ro1 (
   .en(en),
   .out(out[1]),
);

not_3_ro ro2 (
   .en(en),
   .out(out[2]),
);

not_3_ro ro3 (
   .en(en),
   .out(out[3]),
);

not_3_ro ro4 (
   .en(en),
   .out(out[4]),
);

not_3_ro ro5 (
   .en(en),
   .out(out[5]),
);

not_3_ro ro6 (
   .en(en),
   .out(out[6]),
);

not_3_ro ro7 (
   .en(en),
   .out(out[7]),
);

not_3_ro ro8 (
   .en(en),
   .out(out[8]),
);

not_3_ro ro9 (
   .en(en),
   .out(out[9]),
);

not_3_ro ro10 (
   .en(en),
   .out(out[10]),
);

not_3_ro ro11 (
   .en(en),
   .out(out[11]),
);

not_3_ro ro12 (
   .en(en),
   .out(out[12]),
);

not_3_ro ro13 (
   .en(en),
   .out(out[13]),
);

not_3_ro ro14 (
   .en(en),
   .out(out[14]),
);

not_3_ro ro15 (
   .en(en),
   .out(out[15]),
);

not_3_ro ro16 (
   .en(en),
   .out(out[16]),
);

not_3_ro ro17 (
   .en(en),
   .out(out[17]),
);

not_3_ro ro18 (
   .en(en),
   .out(out[18]),
);

not_3_ro ro19 (
   .en(en),
   .out(out[19]),
);

not_3_ro ro20 (
   .en(en),
   .out(out[20]),
);

not_3_ro ro21 (
   .en(en),
   .out(out[21]),
);

not_3_ro ro22 (
   .en(en),
   .out(out[22]),
);

not_3_ro ro23 (
   .en(en),
   .out(out[23]),
);

not_3_ro ro24 (
   .en(en),
   .out(out[24]),
);

not_3_ro ro25 (
   .en(en),
   .out(out[25]),
);

not_3_ro ro26 (
   .en(en),
   .out(out[26]),
);

not_3_ro ro27 (
   .en(en),
   .out(out[27]),
);

not_3_ro ro28 (
   .en(en),
   .out(out[28]),
);

not_3_ro ro29 (
   .en(en),
   .out(out[29]),
);

not_3_ro ro30 (
   .en(en),
   .out(out[30]),
);

not_3_ro ro31 (
   .en(en),
   .out(out[31]),
);

not_3_ro ro32 (
   .en(en),
   .out(out[32]),
);

not_3_ro ro33 (
   .en(en),
   .out(out[33]),
);

not_3_ro ro34 (
   .en(en),
   .out(out[34]),
);

not_3_ro ro35 (
   .en(en),
   .out(out[35]),
);

not_3_ro ro36 (
   .en(en),
   .out(out[36]),
);

not_3_ro ro37 (
   .en(en),
   .out(out[37]),
);

not_3_ro ro38 (
   .en(en),
   .out(out[38]),
);

not_3_ro ro39 (
   .en(en),
   .out(out[39]),
);

not_3_ro ro40 (
   .en(en),
   .out(out[40]),
);

not_3_ro ro41 (
   .en(en),
   .out(out[41]),
);

not_3_ro ro42 (
   .en(en),
   .out(out[42]),
);

not_3_ro ro43 (
   .en(en),
   .out(out[43]),
);

not_3_ro ro44 (
   .en(en),
   .out(out[44]),
);

not_3_ro ro45 (
   .en(en),
   .out(out[45]),
);

not_3_ro ro46 (
   .en(en),
   .out(out[46]),
);

not_3_ro ro47 (
   .en(en),
   .out(out[47]),
);

not_3_ro ro48 (
   .en(en),
   .out(out[48]),
);

not_3_ro ro49 (
   .en(en),
   .out(out[49]),
);

not_3_ro ro50 (
   .en(en),
   .out(out[50]),
);

not_3_ro ro51 (
   .en(en),
   .out(out[51]),
);

not_3_ro ro52 (
   .en(en),
   .out(out[52]),
);

not_3_ro ro53 (
   .en(en),
   .out(out[53]),
);

not_3_ro ro54 (
   .en(en),
   .out(out[54]),
);

not_3_ro ro55 (
   .en(en),
   .out(out[55]),
);

not_3_ro ro56 (
   .en(en),
   .out(out[56]),
);

not_3_ro ro57 (
   .en(en),
   .out(out[57]),
);

not_3_ro ro58 (
   .en(en),
   .out(out[58]),
);

not_3_ro ro59 (
   .en(en),
   .out(out[59]),
);

not_3_ro ro60 (
   .en(en),
   .out(out[60]),
);

not_3_ro ro61 (
   .en(en),
   .out(out[61]),
);

not_3_ro ro62 (
   .en(en),
   .out(out[62]),
);

not_3_ro ro63 (
   .en(en),
   .out(out[63]),
);

not_3_ro ro64 (
   .en(en),
   .out(out[64]),
);

not_3_ro ro65 (
   .en(en),
   .out(out[65]),
);

not_3_ro ro66 (
   .en(en),
   .out(out[66]),
);

not_3_ro ro67 (
   .en(en),
   .out(out[67]),
);

not_3_ro ro68 (
   .en(en),
   .out(out[68]),
);

not_3_ro ro69 (
   .en(en),
   .out(out[69]),
);

not_3_ro ro70 (
   .en(en),
   .out(out[70]),
);

not_3_ro ro71 (
   .en(en),
   .out(out[71]),
);

not_3_ro ro72 (
   .en(en),
   .out(out[72]),
);

not_3_ro ro73 (
   .en(en),
   .out(out[73]),
);

not_3_ro ro74 (
   .en(en),
   .out(out[74]),
);

not_3_ro ro75 (
   .en(en),
   .out(out[75]),
);

not_3_ro ro76 (
   .en(en),
   .out(out[76]),
);

not_3_ro ro77 (
   .en(en),
   .out(out[77]),
);

not_3_ro ro78 (
   .en(en),
   .out(out[78]),
);

not_3_ro ro79 (
   .en(en),
   .out(out[79]),
);

not_3_ro ro80 (
   .en(en),
   .out(out[80]),
);

not_3_ro ro81 (
   .en(en),
   .out(out[81]),
);

not_3_ro ro82 (
   .en(en),
   .out(out[82]),
);

not_3_ro ro83 (
   .en(en),
   .out(out[83]),
);

not_3_ro ro84 (
   .en(en),
   .out(out[84]),
);

not_3_ro ro85 (
   .en(en),
   .out(out[85]),
);

not_3_ro ro86 (
   .en(en),
   .out(out[86]),
);

not_3_ro ro87 (
   .en(en),
   .out(out[87]),
);

not_3_ro ro88 (
   .en(en),
   .out(out[88]),
);

not_3_ro ro89 (
   .en(en),
   .out(out[89]),
);

not_3_ro ro90 (
   .en(en),
   .out(out[90]),
);

not_3_ro ro91 (
   .en(en),
   .out(out[91]),
);

not_3_ro ro92 (
   .en(en),
   .out(out[92]),
);

not_3_ro ro93 (
   .en(en),
   .out(out[93]),
);

not_3_ro ro94 (
   .en(en),
   .out(out[94]),
);

not_3_ro ro95 (
   .en(en),
   .out(out[95]),
);

not_3_ro ro96 (
   .en(en),
   .out(out[96]),
);

not_3_ro ro97 (
   .en(en),
   .out(out[97]),
);

not_3_ro ro98 (
   .en(en),
   .out(out[98]),
);

not_3_ro ro99 (
   .en(en),
   .out(out[99]),
);

not_3_ro ro100 (
   .en(en),
   .out(out[100]),
);

not_3_ro ro101 (
   .en(en),
   .out(out[101]),
);

not_3_ro ro102 (
   .en(en),
   .out(out[102]),
);

not_3_ro ro103 (
   .en(en),
   .out(out[103]),
);

not_3_ro ro104 (
   .en(en),
   .out(out[104]),
);

not_3_ro ro105 (
   .en(en),
   .out(out[105]),
);

not_3_ro ro106 (
   .en(en),
   .out(out[106]),
);

not_3_ro ro107 (
   .en(en),
   .out(out[107]),
);

not_3_ro ro108 (
   .en(en),
   .out(out[108]),
);

not_3_ro ro109 (
   .en(en),
   .out(out[109]),
);

not_3_ro ro110 (
   .en(en),
   .out(out[110]),
);

not_3_ro ro111 (
   .en(en),
   .out(out[111]),
);

not_3_ro ro112 (
   .en(en),
   .out(out[112]),
);

not_3_ro ro113 (
   .en(en),
   .out(out[113]),
);

not_3_ro ro114 (
   .en(en),
   .out(out[114]),
);

not_3_ro ro115 (
   .en(en),
   .out(out[115]),
);

not_3_ro ro116 (
   .en(en),
   .out(out[116]),
);

not_3_ro ro117 (
   .en(en),
   .out(out[117]),
);

not_3_ro ro118 (
   .en(en),
   .out(out[118]),
);

not_3_ro ro119 (
   .en(en),
   .out(out[119]),
);

not_3_ro ro120 (
   .en(en),
   .out(out[120]),
);

not_3_ro ro121 (
   .en(en),
   .out(out[121]),
);

not_3_ro ro122 (
   .en(en),
   .out(out[122]),
);

not_3_ro ro123 (
   .en(en),
   .out(out[123]),
);

not_3_ro ro124 (
   .en(en),
   .out(out[124]),
);

not_3_ro ro125 (
   .en(en),
   .out(out[125]),
);

not_3_ro ro126 (
   .en(en),
   .out(out[126]),
);

not_3_ro ro127 (
   .en(en),
   .out(out[127]),
);

not_3_ro ro128 (
   .en(en),
   .out(out[128]),
);

not_3_ro ro129 (
   .en(en),
   .out(out[129]),
);

not_3_ro ro130 (
   .en(en),
   .out(out[130]),
);

not_3_ro ro131 (
   .en(en),
   .out(out[131]),
);

not_3_ro ro132 (
   .en(en),
   .out(out[132]),
);

not_3_ro ro133 (
   .en(en),
   .out(out[133]),
);

not_3_ro ro134 (
   .en(en),
   .out(out[134]),
);

not_3_ro ro135 (
   .en(en),
   .out(out[135]),
);

not_3_ro ro136 (
   .en(en),
   .out(out[136]),
);

not_3_ro ro137 (
   .en(en),
   .out(out[137]),
);

not_3_ro ro138 (
   .en(en),
   .out(out[138]),
);

not_3_ro ro139 (
   .en(en),
   .out(out[139]),
);

not_3_ro ro140 (
   .en(en),
   .out(out[140]),
);

not_3_ro ro141 (
   .en(en),
   .out(out[141]),
);

not_3_ro ro142 (
   .en(en),
   .out(out[142]),
);

not_3_ro ro143 (
   .en(en),
   .out(out[143]),
);

not_3_ro ro144 (
   .en(en),
   .out(out[144]),
);

not_3_ro ro145 (
   .en(en),
   .out(out[145]),
);

not_3_ro ro146 (
   .en(en),
   .out(out[146]),
);

not_3_ro ro147 (
   .en(en),
   .out(out[147]),
);

not_3_ro ro148 (
   .en(en),
   .out(out[148]),
);

not_3_ro ro149 (
   .en(en),
   .out(out[149]),
);

not_3_ro ro150 (
   .en(en),
   .out(out[150]),
);

not_3_ro ro151 (
   .en(en),
   .out(out[151]),
);

not_3_ro ro152 (
   .en(en),
   .out(out[152]),
);

not_3_ro ro153 (
   .en(en),
   .out(out[153]),
);

not_3_ro ro154 (
   .en(en),
   .out(out[154]),
);

not_3_ro ro155 (
   .en(en),
   .out(out[155]),
);

not_3_ro ro156 (
   .en(en),
   .out(out[156]),
);

not_3_ro ro157 (
   .en(en),
   .out(out[157]),
);

not_3_ro ro158 (
   .en(en),
   .out(out[158]),
);

not_3_ro ro159 (
   .en(en),
   .out(out[159]),
);

not_3_ro ro160 (
   .en(en),
   .out(out[160]),
);

not_3_ro ro161 (
   .en(en),
   .out(out[161]),
);

not_3_ro ro162 (
   .en(en),
   .out(out[162]),
);

not_3_ro ro163 (
   .en(en),
   .out(out[163]),
);

not_3_ro ro164 (
   .en(en),
   .out(out[164]),
);

not_3_ro ro165 (
   .en(en),
   .out(out[165]),
);

not_3_ro ro166 (
   .en(en),
   .out(out[166]),
);

not_3_ro ro167 (
   .en(en),
   .out(out[167]),
);

not_3_ro ro168 (
   .en(en),
   .out(out[168]),
);

not_3_ro ro169 (
   .en(en),
   .out(out[169]),
);

not_3_ro ro170 (
   .en(en),
   .out(out[170]),
);

not_3_ro ro171 (
   .en(en),
   .out(out[171]),
);

not_3_ro ro172 (
   .en(en),
   .out(out[172]),
);

not_3_ro ro173 (
   .en(en),
   .out(out[173]),
);

not_3_ro ro174 (
   .en(en),
   .out(out[174]),
);

not_3_ro ro175 (
   .en(en),
   .out(out[175]),
);

not_3_ro ro176 (
   .en(en),
   .out(out[176]),
);

not_3_ro ro177 (
   .en(en),
   .out(out[177]),
);

not_3_ro ro178 (
   .en(en),
   .out(out[178]),
);

not_3_ro ro179 (
   .en(en),
   .out(out[179]),
);

not_3_ro ro180 (
   .en(en),
   .out(out[180]),
);

not_3_ro ro181 (
   .en(en),
   .out(out[181]),
);

not_3_ro ro182 (
   .en(en),
   .out(out[182]),
);

not_3_ro ro183 (
   .en(en),
   .out(out[183]),
);

not_3_ro ro184 (
   .en(en),
   .out(out[184]),
);

not_3_ro ro185 (
   .en(en),
   .out(out[185]),
);

not_3_ro ro186 (
   .en(en),
   .out(out[186]),
);

not_3_ro ro187 (
   .en(en),
   .out(out[187]),
);

not_3_ro ro188 (
   .en(en),
   .out(out[188]),
);

not_3_ro ro189 (
   .en(en),
   .out(out[189]),
);

assign io_pad[2] = |out;
endmodule
