

module lut_2_ro(
   input en,
   output out,
);

(*keep*)wire connect;
wire test;

assign out = connect;

mux2x0 enable (
   .S(en),
   .A(1'b0),
   .B(connect),
   .Q(test),
);

LUT2 #(
   .INIT(4'b0001)
) ro (
   .I0(test),
   .I1(1'b0),
   .O(connect)
);
endmodule

 
module MODULE_top(
   io_pad
);

// GPIO
inout    wire     [31:0]      io_pad      ;

wire [149:0] out;

// Initialize 48MHz clock
wire                                    CLK        ;
wire                                    CLK_RST    ;

qlal4s3b_cell_macro u_qlal4s3b_cell_macro (
    // FB Clocks
    .Sys_Clk0                  ( CLK                       ), // output
    .Sys_Clk0_Rst              ( CLK_RST                   ), // output
);

reg  [31:0] counter;

reg en;

always @(posedge CLK) begin
   if (counter > 100000000) begin
      en <= 1;
   end
   counter = counter + 1;
end

lut_2_ro ro1(
   .en(en),
   .out(out[0]),
);

lut_2_ro ro2(
   .en(en),
   .out(out[1]),
);

lut_2_ro ro3(
   .en(en),
   .out(out[2]),
);

lut_2_ro ro4(
   .en(en),
   .out(out[3]),
);

lut_2_ro ro5(
   .en(en),
   .out(out[4]),
);

lut_2_ro ro6(
   .en(en),
   .out(out[5]),
);

lut_2_ro ro7(
   .en(en),
   .out(out[6]),
);

lut_2_ro ro8(
   .en(en),
   .out(out[7]),
);

lut_2_ro ro9(
   .en(en),
   .out(out[8]),
);

lut_2_ro ro10(
   .en(en),
   .out(out[9]),
);

lut_2_ro ro11(
   .en(en),
   .out(out[10]),
);

lut_2_ro ro12(
   .en(en),
   .out(out[11]),
);

lut_2_ro ro13(
   .en(en),
   .out(out[12]),
);

lut_2_ro ro14(
   .en(en),
   .out(out[13]),
);

lut_2_ro ro15(
   .en(en),
   .out(out[14]),
);

lut_2_ro ro16(
   .en(en),
   .out(out[15]),
);

lut_2_ro ro17(
   .en(en),
   .out(out[16]),
);

lut_2_ro ro18(
   .en(en),
   .out(out[17]),
);

lut_2_ro ro19(
   .en(en),
   .out(out[18]),
);

lut_2_ro ro20(
   .en(en),
   .out(out[19]),
);

lut_2_ro ro21(
   .en(en),
   .out(out[20]),
);

lut_2_ro ro22(
   .en(en),
   .out(out[21]),
);

lut_2_ro ro23(
   .en(en),
   .out(out[22]),
);

lut_2_ro ro24(
   .en(en),
   .out(out[23]),
);

lut_2_ro ro25(
   .en(en),
   .out(out[24]),
);

lut_2_ro ro26(
   .en(en),
   .out(out[25]),
);

lut_2_ro ro27(
   .en(en),
   .out(out[26]),
);

lut_2_ro ro28(
   .en(en),
   .out(out[27]),
);

lut_2_ro ro29(
   .en(en),
   .out(out[28]),
);

lut_2_ro ro30(
   .en(en),
   .out(out[29]),
);

lut_2_ro ro31(
   .en(en),
   .out(out[30]),
);

lut_2_ro ro32(
   .en(en),
   .out(out[31]),
);

lut_2_ro ro33(
   .en(en),
   .out(out[32]),
);

lut_2_ro ro34(
   .en(en),
   .out(out[33]),
);

lut_2_ro ro35(
   .en(en),
   .out(out[34]),
);

lut_2_ro ro36(
   .en(en),
   .out(out[35]),
);

lut_2_ro ro37(
   .en(en),
   .out(out[36]),
);

lut_2_ro ro38(
   .en(en),
   .out(out[37]),
);

lut_2_ro ro39(
   .en(en),
   .out(out[38]),
);

lut_2_ro ro40(
   .en(en),
   .out(out[39]),
);

lut_2_ro ro41(
   .en(en),
   .out(out[40]),
);

lut_2_ro ro42(
   .en(en),
   .out(out[41]),
);

lut_2_ro ro43(
   .en(en),
   .out(out[42]),
);

lut_2_ro ro44(
   .en(en),
   .out(out[43]),
);

lut_2_ro ro45(
   .en(en),
   .out(out[44]),
);

lut_2_ro ro46(
   .en(en),
   .out(out[45]),
);

lut_2_ro ro47(
   .en(en),
   .out(out[46]),
);

lut_2_ro ro48(
   .en(en),
   .out(out[47]),
);

lut_2_ro ro49(
   .en(en),
   .out(out[48]),
);

lut_2_ro ro50(
   .en(en),
   .out(out[49]),
);

lut_2_ro ro51(
   .en(en),
   .out(out[50]),
);

lut_2_ro ro52(
   .en(en),
   .out(out[51]),
);

lut_2_ro ro53(
   .en(en),
   .out(out[52]),
);

lut_2_ro ro54(
   .en(en),
   .out(out[53]),
);

lut_2_ro ro55(
   .en(en),
   .out(out[54]),
);

lut_2_ro ro56(
   .en(en),
   .out(out[55]),
);

lut_2_ro ro57(
   .en(en),
   .out(out[56]),
);

lut_2_ro ro58(
   .en(en),
   .out(out[57]),
);

lut_2_ro ro59(
   .en(en),
   .out(out[58]),
);

lut_2_ro ro60(
   .en(en),
   .out(out[59]),
);

lut_2_ro ro61(
   .en(en),
   .out(out[60]),
);

lut_2_ro ro62(
   .en(en),
   .out(out[61]),
);

lut_2_ro ro63(
   .en(en),
   .out(out[62]),
);

lut_2_ro ro64(
   .en(en),
   .out(out[63]),
);

lut_2_ro ro65(
   .en(en),
   .out(out[64]),
);

lut_2_ro ro66(
   .en(en),
   .out(out[65]),
);

lut_2_ro ro67(
   .en(en),
   .out(out[66]),
);

lut_2_ro ro68(
   .en(en),
   .out(out[67]),
);

lut_2_ro ro69(
   .en(en),
   .out(out[68]),
);

lut_2_ro ro70(
   .en(en),
   .out(out[69]),
);

lut_2_ro ro71(
   .en(en),
   .out(out[70]),
);

lut_2_ro ro72(
   .en(en),
   .out(out[71]),
);

lut_2_ro ro73(
   .en(en),
   .out(out[72]),
);

lut_2_ro ro74(
   .en(en),
   .out(out[73]),
);

lut_2_ro ro75(
   .en(en),
   .out(out[74]),
);

lut_2_ro ro76(
   .en(en),
   .out(out[75]),
);

lut_2_ro ro77(
   .en(en),
   .out(out[76]),
);

lut_2_ro ro78(
   .en(en),
   .out(out[77]),
);

lut_2_ro ro79(
   .en(en),
   .out(out[78]),
);

lut_2_ro ro80(
   .en(en),
   .out(out[79]),
);

lut_2_ro ro81(
   .en(en),
   .out(out[80]),
);

lut_2_ro ro82(
   .en(en),
   .out(out[81]),
);

lut_2_ro ro83(
   .en(en),
   .out(out[82]),
);

lut_2_ro ro84(
   .en(en),
   .out(out[83]),
);

lut_2_ro ro85(
   .en(en),
   .out(out[84]),
);

lut_2_ro ro86(
   .en(en),
   .out(out[85]),
);

lut_2_ro ro87(
   .en(en),
   .out(out[86]),
);

lut_2_ro ro88(
   .en(en),
   .out(out[87]),
);

lut_2_ro ro89(
   .en(en),
   .out(out[88]),
);

lut_2_ro ro90(
   .en(en),
   .out(out[89]),
);

lut_2_ro ro91(
   .en(en),
   .out(out[90]),
);

lut_2_ro ro92(
   .en(en),
   .out(out[91]),
);

lut_2_ro ro93(
   .en(en),
   .out(out[92]),
);

lut_2_ro ro94(
   .en(en),
   .out(out[93]),
);

lut_2_ro ro95(
   .en(en),
   .out(out[94]),
);

lut_2_ro ro96(
   .en(en),
   .out(out[95]),
);

lut_2_ro ro97(
   .en(en),
   .out(out[96]),
);

lut_2_ro ro98(
   .en(en),
   .out(out[97]),
);

lut_2_ro ro99(
   .en(en),
   .out(out[98]),
);

lut_2_ro ro100(
   .en(en),
   .out(out[99]),
);

lut_2_ro ro101(
   .en(en),
   .out(out[100]),
);

lut_2_ro ro102(
   .en(en),
   .out(out[101]),
);

lut_2_ro ro103(
   .en(en),
   .out(out[102]),
);

lut_2_ro ro104(
   .en(en),
   .out(out[103]),
);

lut_2_ro ro105(
   .en(en),
   .out(out[104]),
);

lut_2_ro ro106(
   .en(en),
   .out(out[105]),
);

lut_2_ro ro107(
   .en(en),
   .out(out[106]),
);

lut_2_ro ro108(
   .en(en),
   .out(out[107]),
);

lut_2_ro ro109(
   .en(en),
   .out(out[108]),
);

lut_2_ro ro110(
   .en(en),
   .out(out[109]),
);

lut_2_ro ro111(
   .en(en),
   .out(out[110]),
);

lut_2_ro ro112(
   .en(en),
   .out(out[111]),
);

lut_2_ro ro113(
   .en(en),
   .out(out[112]),
);

lut_2_ro ro114(
   .en(en),
   .out(out[113]),
);

lut_2_ro ro115(
   .en(en),
   .out(out[114]),
);

lut_2_ro ro116(
   .en(en),
   .out(out[115]),
);

lut_2_ro ro117(
   .en(en),
   .out(out[116]),
);

lut_2_ro ro118(
   .en(en),
   .out(out[117]),
);

lut_2_ro ro119(
   .en(en),
   .out(out[118]),
);

lut_2_ro ro120(
   .en(en),
   .out(out[119]),
);

lut_2_ro ro121(
   .en(en),
   .out(out[120]),
);

lut_2_ro ro122(
   .en(en),
   .out(out[121]),
);

lut_2_ro ro123(
   .en(en),
   .out(out[122]),
);

lut_2_ro ro124(
   .en(en),
   .out(out[123]),
);

lut_2_ro ro125(
   .en(en),
   .out(out[124]),
);

lut_2_ro ro126(
   .en(en),
   .out(out[125]),
);

lut_2_ro ro127(
   .en(en),
   .out(out[126]),
);

lut_2_ro ro128(
   .en(en),
   .out(out[127]),
);

lut_2_ro ro129(
   .en(en),
   .out(out[128]),
);

lut_2_ro ro130(
   .en(en),
   .out(out[129]),
);

lut_2_ro ro131(
   .en(en),
   .out(out[130]),
);

lut_2_ro ro132(
   .en(en),
   .out(out[131]),
);

lut_2_ro ro133(
   .en(en),
   .out(out[132]),
);

lut_2_ro ro134(
   .en(en),
   .out(out[133]),
);

lut_2_ro ro135(
   .en(en),
   .out(out[134]),
);

lut_2_ro ro136(
   .en(en),
   .out(out[135]),
);

lut_2_ro ro137(
   .en(en),
   .out(out[136]),
);

lut_2_ro ro138(
   .en(en),
   .out(out[137]),
);

lut_2_ro ro139(
   .en(en),
   .out(out[138]),
);

lut_2_ro ro140(
   .en(en),
   .out(out[139]),
);

lut_2_ro ro141(
   .en(en),
   .out(out[140]),
);

lut_2_ro ro142(
   .en(en),
   .out(out[141]),
);

lut_2_ro ro143(
   .en(en),
   .out(out[142]),
);

lut_2_ro ro144(
   .en(en),
   .out(out[143]),
);

lut_2_ro ro145(
   .en(en),
   .out(out[144]),
);

lut_2_ro ro146(
   .en(en),
   .out(out[145]),
);

lut_2_ro ro147(
   .en(en),
   .out(out[146]),
);

lut_2_ro ro148(
   .en(en),
   .out(out[147]),
);

lut_2_ro ro149(
   .en(en),
   .out(out[148]),
);

lut_2_ro ro150(
   .en(en),
   .out(out[149]),
);
assign io_pad[13] = |out;
endmodule
